
module s15850 ( CK, g100, g101, g102, g103, g10377, g10379, g104, g10455, 
        g10457, g10459, g10461, g10463, g10465, g10628, g10801, g109, g11163, 
        g11206, g11489, g1170, g1173, g1176, g1179, g1182, g1185, g1188, g1191, 
        g1194, g1197, g1200, g1203, g1696, g1700, g1712, g18, g1957, g1960, 
        g1961, g23, g2355, g2601, g2602, g2603, g2604, g2605, g2606, g2607, 
        g2608, g2609, g2610, g2611, g2612, g2648, g27, g28, g29, g2986, g30, 
        g3007, g3069, g31, g3327, g41, g4171, g4172, g4173, g4174, g4175, 
        g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194, 
        g4195, g4196, g4197, g4198, g4199, g42, g4200, g4201, g4202, g4203, 
        g4204, g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, 
        g4214, g4215, g4216, g43, g44, g45, g46, g47, g48, g4887, g4888, g5101, 
        g5105, g5658, g5659, g5816, g6253, g6254, g6255, g6256, g6257, g6258, 
        g6259, g6260, g6261, g6262, g6263, g6264, g6265, g6266, g6267, g6268, 
        g6269, g6270, g6271, g6272, g6273, g6274, g6275, g6276, g6277, g6278, 
        g6279, g6280, g6281, g6282, g6283, g6284, g6285, g6842, g6920, g6926, 
        g6932, g6942, g6949, g6955, g741, g742, g743, g744, g750, g7744, g8061, 
        g8062, g82, g8271, g83, g8313, g8316, g8318, g8323, g8328, g8331, 
        g8335, g8340, g8347, g8349, g8352, g84, g85, g8561, g8562, g8563, 
        g8564, g8565, g8566, g86, g87, g872, g873, g877, g88, g881, g886, g889, 
        g89, g892, g895, g8976, g8977, g8978, g8979, g898, g8980, g8981, g8982, 
        g8983, g8984, g8985, g8986, g90, g901, g904, g907, g91, g910, g913, 
        g916, g919, g92, g922, g925, g93, g94, g9451, g95, g96, g99, g9961, 
        test_se, test_si1, test_so1, test_si2, test_so2, test_si3, test_so3, 
        test_si4, test_so4, test_si5, test_so5, test_si6, test_so6, test_si7, 
        test_so7, test_si8, test_so8, test_si9, test_so9, test_si10, test_so10
 );
  input CK, g100, g101, g102, g103, g104, g109, g1170, g1173, g1176, g1179,
         g1182, g1185, g1188, g1191, g1194, g1197, g1200, g1203, g1696, g1700,
         g1712, g18, g1960, g1961, g23, g27, g28, g29, g30, g31, g41, g42, g43,
         g44, g45, g46, g47, g48, g741, g742, g743, g744, g750, g82, g83, g84,
         g85, g86, g87, g872, g873, g877, g88, g881, g886, g889, g89, g892,
         g895, g898, g90, g901, g904, g907, g91, g910, g913, g916, g919, g92,
         g922, g925, g93, g94, g95, g96, g99, test_se, test_si1, test_si2,
         test_si3, test_si4, test_si5, test_si6, test_si7, test_si8, test_si9,
         test_si10;
  output g10377, g10379, g10455, g10457, g10459, g10461, g10463, g10465,
         g10628, g10801, g11163, g11206, g11489, g1957, g2355, g2601, g2602,
         g2603, g2604, g2605, g2606, g2607, g2608, g2609, g2610, g2611, g2612,
         g2648, g2986, g3007, g3069, g3327, g4171, g4172, g4173, g4174, g4175,
         g4176, g4177, g4178, g4179, g4180, g4181, g4191, g4192, g4193, g4194,
         g4195, g4196, g4197, g4198, g4199, g4200, g4201, g4202, g4203, g4204,
         g4205, g4206, g4207, g4208, g4209, g4210, g4211, g4212, g4213, g4214,
         g4215, g4216, g4887, g4888, g5101, g5105, g5658, g5659, g5816, g6253,
         g6254, g6255, g6256, g6257, g6258, g6259, g6260, g6261, g6262, g6263,
         g6264, g6265, g6266, g6267, g6268, g6269, g6270, g6271, g6272, g6273,
         g6274, g6275, g6276, g6277, g6278, g6279, g6280, g6281, g6282, g6283,
         g6284, g6285, g6842, g6920, g6926, g6932, g6942, g6949, g6955, g7744,
         g8061, g8062, g8271, g8313, g8316, g8318, g8323, g8328, g8331, g8335,
         g8340, g8347, g8349, g8352, g8561, g8562, g8563, g8564, g8565, g8566,
         g8976, g8977, g8978, g8979, g8980, g8981, g8982, g8983, g8984, g8985,
         g8986, g9451, g9961, test_so1, test_so2, test_so3, test_so4, test_so5,
         test_so6, test_so7, test_so8, test_so9, test_so10;
  wire   N599, g1289, g1882, g312, g452, g11257, g123, g207, g713, g1153,
         g1744, g1558, g695, g461, g940, g976, g709, g8432, g1092, g1574,
         g1864, g369, g1580, g1736, g1424, g1737, g1672, g1077, g1231, g4,
         g1104, g1304, g7290, g243, g1499, g1444, g1543, g315, g1534, g622,
         g1927, g1660, g278, g1436, g718, g8433, g554, g496, g11333, g981,
         g829, g1095, g704, g1265, g7302, g1786, g682, g8429, g1296, g7292,
         g327, g1389, g1371, g1956, g1955, g1675, g354, g113, g639, g1684,
         g1639, g1791, g248, g1707, g1759, g351, g1604, g1098, g932, g1896,
         g8282, g736, g8435, g1019, g745, g1419, g32, g1086, g1486, g1730,
         g1504, g1470, g822, g1678, g174, g1766, g1801, g186, g959, g1407,
         g1868, g1718, g396, g11265, g1015, g1415, g1227, g1721, g284, g426,
         g11256, g219, g1360, g806, g1428, g1564, g1741, g225, g281, g1308,
         g611, g1217, g1589, g1466, g1571, g1861, g1448, g1133, g1333, g153,
         g962, g486, g11331, g471, g1397, g1950, g8288, g756, g755, g1101,
         g549, g105, g1669, g1531, g1458, g572, g1011, g1411, g1074, g444,
         g11259, g1474, g1080, g1713, g333, g269, g401, g11266, g1857, g9,
         g664, g965, g1400, g309, g814, g231, g557, g869, g875, g1383, g158,
         g627, g1023, g259, g1327, g654, g293, g1346, g1633, g1753, g1508,
         g1240, g7297, g538, g11326, g416, g11269, g542, g11325, g1681, g374,
         g563, g1914, g8284, g530, g11328, g575, g1936, g1317, g1356, g357,
         g386, g11263, g1601, g166, g501, g11334, g262, g1840, g318, g794,
         g302, g342, g1250, g7299, g1163, g1032, g1432, g1453, g363, g330,
         g1157, g928, g261, g516, g11337, g254, g861, g1627, g1292, g7293,
         g290, g1583, g466, g1561, g1546, g287, g560, g617, g336, g456, g305,
         g345, g8, g255, g1945, g1738, g1478, g1690, g1482, g1110, g296, g1663,
         g700, g8431, g1762, g360, g192, g1657, g722, g566, g1089, g1071, g986,
         g971, g143, g1814, g1212, g1918, g1822, g237, g746, g1462, g178, g366,
         g837, g599, g1854, g944, g1941, g8287, g170, g1520, g686, g953, g1958,
         g1765, g1733, g7303, g1610, g1796, g1324, g1540, g491, g11332, g213,
         g1781, g1900, g1245, g7298, g148, g833, g1923, g8285, g936, g1314,
         g849, g1336, g272, g1806, g826, g1887, g8281, g968, g1137, g1891,
         g1255, g7300, g257, g874, g591, g731, g636, g1218, g605, g182, g950,
         g1129, g857, g448, g11258, g1828, g1727, g1592, g1703, g1932, g8286,
         g1624, g440, g11260, g476, g11338, g119, g668, g139, g1149, g263,
         g818, g1747, g802, g275, g1524, g1577, g810, g391, g11264, g658,
         g1386, g253, g1125, g201, g1280, g7295, g1083, g650, g1636, g853,
         g421, g11270, g956, g378, g1756, g841, g1027, g1003, g1403, g1145,
         g1107, g1223, g406, g11267, g1811, g1654, g197, g1595, g1537, g727,
         g8434, g798, g481, g11324, g1330, g845, g1512, g1490, g1166, g348,
         g1260, g7301, g260, g131, g258, g521, g11330, g1318, g1872, g677,
         g1549, g947, g1834, g1598, g1121, g1321, g506, g11335, g546, g1909,
         g1552, g1687, g1586, g324, g1141, g1341, g1710, g135, g525, g11329,
         g1607, g321, g1275, g11443, g1615, g382, g266, g1284, g7294, g673,
         g8428, g162, g411, g11268, g431, g11262, g1905, g8283, g1515, g1630,
         g991, g1300, g7291, g339, g256, g1750, g1440, g1666, g1528, g1351,
         g127, g1618, g1235, g7296, g299, g435, g11261, g1555, g995, g1621,
         g643, g1494, g1567, g691, g8430, g534, g11327, g1776, g569, g1160, g1,
         g511, g11336, g1724, g12, g1878, g4500, g5529, g4338, g8147, g6551,
         g10865, g8054, g7709, g4940, g6481, g6529, g10707, g6949, g8940,
         g10855, g6920, g6907, g6155, g6638, g11647, g6910, g6828, g10800,
         g8019, g6821, g11478, g6516, g8244, g8631, g10793, g5910, g2478,
         g10726, g6824, g9961, g6759, g6502, g10797, g4471, g10780, g11625,
         g11372, g10771, g11293, g8173, g6533, g8245, g10767, g6000, g4490,
         g4903, g10720, g6934, g6123, g6838, g4905, g10798, g10785, g7204,
         g6830, g8944, g5543, g8921, g6096, g6942, g6733, g6823, g4890, g3381,
         g10863, g8039, g6526, g10664, g7189, g8923, g5173, g4264, g6755,
         g11514, g4506, g4465, g6902, g6015, g11340, g6542, g6507, g5556,
         g8505, g11641, g10765, g11305, g6126, g8060, g7191, g6469, g4498,
         g6627, g4893, g5194, g6901, g8043, g6929, g8049, g6786, g6234, g10864,
         g8984, g10862, g10721, g8051, g6541, g10773, g8193, g6523, g5404,
         g11393, g4334, g6908, g8768, g8885, g6333, g6045, g7590, g6468,
         g10782, g6672, g6840, g5914, g7705, g6038, g6471, g11303, g10663,
         g8920, g4283, g4484, g5396, g8045, g7843, g6932, g6537, g4902, g6080,
         g6059, g4089, g5126, g10866, g11603, g6332, g4231, g11488, g6955,
         g5918, g6894, g4076, g6534, g6928, g6926, g8055, g11291, g6833, g6918,
         g6915, g6911, g7441, g5996, g8047, g6653, g6832, g11481, g6478, g6897,
         g6042, g4342, g4330, g11609, g10859, g6054, g6508, g6531, g8050,
         g11376, g8559, g7032, g4293, g5390, g8767, g4480, g11483, g5392,
         g10776, g6513, g9272, g10898, g8052, g4325, g8766, g6205, g8820,
         g9124, g6839, g6522, g10936, g11320, g6841, g8769, g6224, g11349,
         g6470, g5755, g6515, g10791, g7632, g11485, g6331, g8053, g5763,
         g6480, g6795, g8194, g8938, g4238, g8775, g4891, g11290, g6501, g6334,
         g10719, g4274, g8765, g6916, g11308, g10784, g6820, g4340, g6922,
         g6747, g11391, g8649, g9555, g6071, g10858, g8926, g4239, g11602,
         g8041, g8922, g5536, g11605, g8048, g6528, g6524, g7219, g8046,
         g11482, g4477, g6923, g4255, g8937, g6538, g11306, g7183, g6895,
         g6179, g9721, g8776, g6827, g4309, g7244, g7586, g7930, g11300,
         g10718, g5445, g6088, g6679, g11636, g9266, g11608, g8059, g8771,
         g6035, g6198, g8973, g6834, g5148, g7134, g10795, g10770, g8773,
         g3462, g7143, g8939, g8772, g6093, g6500, g8777, g6244, g11640,
         g11487, g9110, g11380, g9269, g11314, g9150, g11298, g7202, g6819,
         g6243, g6514, g6983, g4473, g8040, g6900, g8042, g6546, g5770, g8889,
         g10711, g11312, g6479, g5849, g6656, g6906, g10717, g8770, g6392,
         g6621, g11610, g11604, g11486, g7581, g10799, g6439, g7133, g8044,
         g8254, g11607, g6193, g4904, g11292, g6822, g6912, g6898, g5421,
         g6924, g11310, g11294, g6026, g8024, g8945, g6525, g5083, g7541,
         g10860, g11579, g11639, g6826, g7626, g6829, g7660, g10722, g8887,
         g11484, g6002, g11606, g6757, g6216, g8941, g4892, g6930, g8250,
         g6049, g8943, g10861, g8779, g6180, g8774, g8260, g6099, g6831, g6068,
         g7137, g6545, g7257, g6909, g8384, g11392, g6506, g8883, g6728,
         g10724, g4556, DFF_121_n1, DFF_122_n1, DFF_126_n1, DFF_136_n1,
         DFF_157_n1, DFF_168_n1, DFF_194_n1, DFF_228_n1, g8271, DFF_242_n1,
         DFF_275_n1, DFF_311_n1, DFF_319_n1, DFF_330_n1, DFF_336_n1,
         DFF_350_n1, DFF_384_n1, DFF_385_n1, DFF_436_n1, DFF_441_n1,
         DFF_445_n1, DFF_452_n1, DFF_489_n1, n517, n518, n519, n520, n521,
         n522, n524, n526, n527, n528, n529, n530, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n542, n544, n545, n546, n547, n548,
         n549, n550, n551, n552, n553, n554, n555, n556, n557, n560, n561,
         n562, n563, n564, n565, n566, n567, n568, n569, n572, n573, n574,
         n575, n576, n577, n578, n579, n580, n581, n583, n592, n594, n595,
         n596, n597, n598, n599, n600, n602, n603, n604, n605, n606, n607,
         n609, n610, n611, n612, n614, n616, n617, n619, n620, n621, n622,
         n623, n624, n625, n627, n629, n630, n631, n632, n633, n634, n643,
         n644, n645, n646, n647, n648, n649, n650, n651, n661, n662, n665,
         n667, n668, n674, n675, n685, n687, n711, n712, n713, n715, n717,
         n718, n719, n720, n721, n725, n744, n793, n794, n795, n796, n797,
         n798, n799, n800, n801, n802, n803, n804, n805, n806, n807, n808,
         n809, n810, n811, n812, n813, n814, n815, n816, n817, n818, n819,
         n820, n821, n822, n823, n824, n825, n826, n827, n828, n829, n830,
         n831, n832, n833, n834, n835, n836, n837, n838, n839, n840, n841,
         n842, n843, n844, n845, n846, n847, n848, n849, n850, n851, n852,
         n853, n854, n855, n856, n857, n858, n859, n860, n861, n862, n863,
         n864, n865, n866, n867, n868, n869, n870, n871, n872, n873, n874,
         n875, n876, n877, n878, n879, n880, n881, n882, n883, n884, n885,
         n886, n887, n888, n889, n890, n891, n892, n893, n894, n895, n896,
         n897, n898, n899, n900, n901, n902, n903, n904, n905, n906, n907,
         n908, n909, n910, n911, n912, n913, n914, n915, n916, n917, n918,
         n919, n920, n921, n922, n923, n924, n925, n926, n927, n928, n929,
         n930, n931, n932, n933, n934, n935, n936, n937, n938, n939, n940,
         n941, n942, n943, n944, n945, n946, n947, n948, n949, n950, n951,
         n952, n953, n954, n955, n956, n957, n958, n959, n960, n961, n962,
         n963, n964, n965, n966, n967, n968, n969, n970, n971, n972, n973,
         n974, n975, n976, n977, n978, n979, n980, n981, n982, n983, n984,
         n985, n986, n987, n988, n989, n990, n991, n992, n993, n994, n995,
         n996, n997, n998, n999, n1000, n1001, n1002, n1003, n1004, n1005,
         n1006, n1007, n1008, n1009, n1010, n1011, n1012, n1013, n1014, n1015,
         n1016, n1017, n1018, n1019, n1020, n1021, n1022, n1023, n1024, n1025,
         n1026, n1027, n1028, n1029, n1030, n1031, n1032, n1033, n1034, n1035,
         n1036, n1037, n1038, n1039, n1040, n1041, n1042, n1043, n1044, n1045,
         n1046, n1047, n1048, n1049, n1050, n1051, n1052, n1053, n1054, n1055,
         n1056, n1057, n1058, n1059, n1060, n1061, n1062, n1063, n1064, n1065,
         n1066, n1067, n1068, n1069, n1070, n1071, n1072, n1073, n1074, n1075,
         n1076, n1077, n1078, n1079, n1080, n1081, n1082, n1083, n1084, n1085,
         n1086, n1087, n1088, n1089, n1090, n1091, n1092, n1093, n1094, n1095,
         n1096, n1097, n1098, n1099, n1100, n1101, n1102, n1103, n1104, n1105,
         n1106, n1107, n1108, n1109, n1110, n1111, n1112, n1113, n1114, n1115,
         n1116, n1117, n1118, n1119, n1120, n1122, n1123, n1124, n1125, n1126,
         n1127, n1128, n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136,
         n1137, n1138, n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146,
         n1147, n1148, n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156,
         n1157, n1158, n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166,
         n1167, n1168, n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176,
         n1177, n1178, n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186,
         n1187, n1188, n1189, n1190, n1191, n1192, n1193, n1195, n1196, n1197,
         n1198, n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207,
         n1208, n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217,
         n1218, n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227,
         n1228, n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237,
         n1238, n1239, n1240, n1241, n1243, n1244, n1245, n1246, n1247, n1248,
         n1249, n1250, n1251, n1252, n1253, n1254, n1255, n1256, n1257, n1258,
         n1259, n1260, n1261, n1262, n1263, n1264, n1265, n1266, n1267, n1268,
         n1269, n1270, n1271, n1272, n1273, n1274, n1275, n1276, n1277, n1278,
         n1279, n1280, n1281, n1282, n1283, n1284, n1285, n1286, n1287, n1288,
         n1289, n1290, n1291, n1292, n1293, n1294, n1295, n1296, n1297, n1298,
         n1299, n1300, n1301, n1302, n1303, n1304, n1305, n1306, n1307, n1308,
         n1309, n1310, n1311, n1312, n1313, n1314, n1315, n1316, n1317, n1318,
         n1319, n1320, n1321, n1322, n1323, n1324, n1325, n1326, n1328, n1329,
         n1330, n1331, n1332, n1333, n1334, n1335, n1336, n1337, n1338, n1339,
         n1340, n1341, n1342, n1343, n1344, n1345, n1346, n1347, n1348, n1349,
         n1350, n1351, n1352, n1353, n1354, n1355, n1356, n1357, n1358, n1359,
         n1360, n1361, n1362, n1363, n1364, n1365, n1366, n1367, n1368, n1369,
         n1370, n1371, n1372, n1373, n1374, n1375, n1376, n1377, n1378, n1379,
         n1380, n1381, n1382, n1383, n1384, n1385, n1386, n1387, n1388, n1389,
         n1390, n1391, n1392, n1393, n1394, n1395, n1396, n1397, n1398, n1399,
         n1402, n1403, n1404, n1405, n1406, n1407, n1408, n1409, n1410, n1411,
         n1412, n1413, n1414, n1415, n1416, n1417, n1418, n1419, n1420, n1421,
         n1422, n1423, n1424, n1425, n1426, n1427, n1428, n1429, n1430, n1431,
         n1432, n1433, n1434, n1436, n1437, n1438, n1439, n1440, n1441, n1442,
         n1443, n1444, n1445, n1446, n1447, n1448, n1449, n1450, n1451, n1452,
         n1453, n1454, n1455, n1459, n1461, n1462, n1463, n1464, n1465, n1466,
         n1467, n1468, n1469, n1470, n1471, n1472, n1473, n1474, n1475, n1476,
         n1477, n1478, n1479, n1480, n1481, n1482, n1483, n1484, n1485, n1486,
         n1487, n1488, n1489, n1490, n1491, n1492, n1493, n1494, n1495, n1496,
         n1497, n1498, n1499, n1500, n1501, n1502, n1503, n1504, n1505, n1506,
         n1507, n1508, n1509, n1510, n1511, n1512, n1513, n1514, n1515, n1516,
         n1517, n1518, n1519, n1520, n1521, n1522, n1523, n1524, n1525, n1526,
         n1527, n1528, n1529, n1530, n1531, n1532, n1533, n1534, n1535, n1536,
         n1537, n1538, n1539, n1540, n1541, n1542, n1543, n1544, n1545, n1546,
         n1547, n1548, n1549, n1550, n1551, n1552, n1553, n1554, n1555, n1556,
         n1557, n1558, n1559, n1560, n1561, n1562, n1563, n1564, n1565, n1566,
         n1567, n1568, n1569, n1570, n1571, n1572, n1573, n1574, n1575, n1576,
         n1577, n1578, n1579, n1580, n1581, n1583, n1585, n1586, n1587, n1588,
         n1590, n1591, n1592, n1593, n1594, n1595, n1596, n1597, n1598, n1599,
         n1600, n1601, n1602, n1603, n1604, n1605, n1606, n1607, n1608, n1609,
         n1610, n1611, n1612, n1613, n1614, n1615, n1616, n1617, n1618, n1619,
         n1620, n1621, n1622, n1623, n1624, n1625, n1626, n1627, n1628, n1629,
         n1630, n1631, n1632, n1633, n1634, n1635, n1636, n1637, n1638, n1639,
         n1640, n1641, n1642, n1643, n1644, n1645, n1646, n1647, n1648, n1649,
         n1650, n1651, n1652, n1653, n1654, n1655, n1656, n1657, n1658, n1659,
         n1660, n1661, n1662, n1663, n1664, n1665, n1666, n1667, n1668, n1669,
         n1670, n1671, n1672, n1673, n1674, n1675, n1676, n1677, n1678, n1679,
         n1680, n1681, n1682, n1683, n1684, n1685, n1686, n1687, n1688, n1689,
         n1690, n1691, n1692, n1693, n1694, n1695, n1696, n1697, n1698, n1699,
         n1700, n1701, n1702, n1703, n1704, n1705, n1706, n1707, n1708, n1709,
         n1710, n1711, n1712, n1713, n1714, n1715, n1716, n1717, n1718, n1719,
         n1720, n1721, n1722, n1723, n1724, n1725, n1727, n1729, n1731, n1733,
         n1735, n1737, n1739, n1741, n1743, n1745, n1747, n1749, n1751, n1753,
         n1755, n1757, n1759, n1761, n1763, n1765, n1767, n1769, n1771, n1773,
         n1775, n1777, n1779, n1781, n1783, n1785, n1787, n1789, n1791, n1793,
         n1795, n1797, n1799, n1801, n1803, n1805, n1807, n1809, n1811, n1813,
         n1815, n1817, n1819, n1821, n1823, n1825, n1827, n1829, n1831, n1833,
         n1835, n1837, g5105, n1839, g5101, n1841, n1843, n1845, n1847, n1849,
         n1851, n1853, n1854, n1855, n1856, n1857, n1858, n1859, n1860, n1861,
         n1862, n1863, n1864, n1865, n1866, n1867, n1868, n1869, n1870, n1871,
         n1872, n1873, n1874, n1875, n1876, n1877, n1878, n1880, n1881, n1882,
         n1883, n1884, n1885, n1886, n1887, n1888, n1889, n1890, n1891, n1892,
         n1893, n1894, n1895, n1896, n1897, n1898, n1899, n1900, n1901, n1902,
         n1903, n1904, n1905, n1906, n1907, n1908, n1909, n1910, n1911, n1912,
         n1913, n1914, n1915, n1916, n1917, n1918, n1919, n1920, n1921, n1922,
         n1923, n1924, n1925, n1926, n1927, n1928, n1929, n1930, n1931, n1932,
         n1933, n1934, n1935, n1936, n1937, n1938, n1939, n1940, n1941, n1942,
         n1943, n1944, n1945, n1946, n1947, n1948, n1949, n1950, n1951, n1952,
         n1953, n1954, n1955, n1956, n1957, n1958, n1959, n1960, n1961, n1962,
         n1963, n1964, n1965, n1966, n1967, n1968, n1969, n1970, n1971, n1972,
         n1973, n1974, n1975, n1976, n1977, n1978, n1979, n1980, n1981, n1982,
         n1983, n1984, n1985, n1986, n1987, n1988, n3016, n3017, n3018, n3019,
         n3020, n3022, n3023, n3024, n3025, n3026, n3027, n3029, n3030, n3031,
         n3033, n3034, n3035, n3036, n3037, n3038, n3040, n3041, n3042, n3044,
         n3045, n3046, n3047, n3048, n3050, n3051, n3053, n3054, n3055, n3056,
         n3057, n3058, n3059, n3061, n3062, n3064, n3065;
  assign g8565 = g6949;
  assign g8561 = g6920;
  assign g9451 = g9961;
  assign g8564 = g6942;
  assign test_so10 = g8984;
  assign g8563 = g6932;
  assign g8566 = g6955;
  assign g8562 = g6926;
  assign g5816 = g8271;
  assign g11489 = 1'b0;
  assign g8062 = g5105;
  assign g8061 = g5101;

  LSDNENX1 U1550 ( .D(g10722), .ENB(n1887), .Q(g10461) );
  LSDNENX1 U1551 ( .D(g10664), .ENB(n1886), .Q(g10379) );
  SDFFX1 DFF_0_Q_reg ( .D(g4556), .SI(test_si1), .SE(test_se), .CLK(CK), .Q(
        g1289), .QN() );
  SDFFX1 DFF_1_Q_reg ( .D(g8943), .SI(g1289), .SE(test_se), .CLK(CK), .Q(g1882), .QN(n1663) );
  SDFFX1 DFF_2_Q_reg ( .D(g255), .SI(g1882), .SE(test_se), .CLK(CK), .Q(g312), 
        .QN() );
  SDFFX1 DFF_3_Q_reg ( .D(g11257), .SI(g312), .SE(test_se), .CLK(CK), .Q(g452), 
        .QN() );
  SDFFX1 DFF_4_Q_reg ( .D(g7032), .SI(g452), .SE(test_se), .CLK(CK), .Q(g123), 
        .QN() );
  SDFFX1 DFF_5_Q_reg ( .D(g6830), .SI(g123), .SE(test_se), .CLK(CK), .Q(g207), 
        .QN() );
  SDFFX1 DFF_6_Q_reg ( .D(g8920), .SI(g207), .SE(test_se), .CLK(CK), .Q(g713), 
        .QN() );
  SDFFX1 DFF_7_Q_reg ( .D(g4340), .SI(g713), .SE(test_se), .CLK(CK), .Q(g1153), 
        .QN(n1686) );
  SDFFX1 DFF_9_Q_reg ( .D(g4239), .SI(g1153), .SE(test_se), .CLK(CK), .Q(g1744), .QN() );
  SDFFX1 DFF_10_Q_reg ( .D(g6538), .SI(g1744), .SE(test_se), .CLK(CK), .Q(
        g1558), .QN() );
  SDFFX1 DFF_11_Q_reg ( .D(g8887), .SI(g1558), .SE(test_se), .CLK(CK), .Q(g695), .QN() );
  SDFFX1 DFF_12_Q_reg ( .D(g11372), .SI(g695), .SE(test_se), .CLK(CK), .Q(g461), .QN(n1594) );
  SDFFX1 DFF_13_Q_reg ( .D(g8260), .SI(g461), .SE(test_se), .CLK(CK), .Q(g940), 
        .QN(n1712) );
  SDFFX1 DFF_14_Q_reg ( .D(g11391), .SI(g940), .SE(test_se), .CLK(CK), .Q(g976), .QN() );
  SDFFX1 DFF_15_Q_reg ( .D(g8432), .SI(g976), .SE(test_se), .CLK(CK), .Q(g709), 
        .QN(n1719) );
  SDFFX1 DFF_16_Q_reg ( .D(g6088), .SI(g709), .SE(test_se), .CLK(CK), .Q(g1092), .QN() );
  SDFFX1 DFF_17_Q_reg ( .D(g6478), .SI(g1092), .SE(test_se), .CLK(CK), .Q(
        g1574), .QN() );
  SDFFX1 DFF_18_Q_reg ( .D(g6795), .SI(g1574), .SE(test_se), .CLK(CK), .Q(
        g1864), .QN() );
  SDFFX1 DFF_19_Q_reg ( .D(g11320), .SI(g1864), .SE(test_se), .CLK(CK), .Q(
        g369), .QN() );
  SDFFX1 DFF_20_Q_reg ( .D(g6500), .SI(g369), .SE(test_se), .CLK(CK), .Q(g1580), .QN() );
  SDFFX1 DFF_21_Q_reg ( .D(g5392), .SI(g1580), .SE(test_se), .CLK(CK), .Q(
        g1736), .QN() );
  SDFFX1 DFF_22_Q_reg ( .D(g10663), .SI(g1736), .SE(test_se), .CLK(CK), .Q(
        n1637), .QN() );
  SDFFX1 DFF_23_Q_reg ( .D(g10782), .SI(n1637), .SE(test_se), .CLK(CK), .Q(
        n3065), .QN(n1590) );
  SDFFX1 DFF_24_Q_reg ( .D(g6216), .SI(n3065), .SE(test_se), .CLK(CK), .Q(
        g1424), .QN() );
  SDFFX1 DFF_25_Q_reg ( .D(g1736), .SI(g1424), .SE(test_se), .CLK(CK), .Q(
        g1737), .QN() );
  SDFFX1 DFF_26_Q_reg ( .D(g10858), .SI(g1737), .SE(test_se), .CLK(CK), .Q(
        g1672), .QN() );
  SDFFX1 DFF_27_Q_reg ( .D(g5914), .SI(g1672), .SE(test_se), .CLK(CK), .Q(
        g1077), .QN() );
  SDFFX1 DFF_28_Q_reg ( .D(g7590), .SI(g1077), .SE(test_se), .CLK(CK), .Q(
        g1231), .QN() );
  SDFFX1 DFF_29_Q_reg ( .D(g6656), .SI(g1231), .SE(test_se), .CLK(CK), .Q(g4), 
        .QN() );
  SDFFX1 DFF_30_Q_reg ( .D(g6728), .SI(g4), .SE(test_se), .CLK(CK), .Q(g4177), 
        .QN() );
  SDFFX1 DFF_31_Q_reg ( .D(g5126), .SI(g4177), .SE(test_se), .CLK(CK), .Q(
        g1104), .QN(n1658) );
  SDFFX1 DFF_32_Q_reg ( .D(g7290), .SI(g1104), .SE(test_se), .CLK(CK), .Q(
        g1304), .QN() );
  SDFFX1 DFF_33_Q_reg ( .D(g6841), .SI(g1304), .SE(test_se), .CLK(CK), .Q(g243), .QN() );
  SDFFX1 DFF_34_Q_reg ( .D(g8041), .SI(g243), .SE(test_se), .CLK(CK), .Q(g1499), .QN() );
  SDFFX1 DFF_36_Q_reg ( .D(g8766), .SI(g1499), .SE(test_se), .CLK(CK), .Q(
        g1444), .QN() );
  SDFFX1 DFF_37_Q_reg ( .D(n524), .SI(g1444), .SE(test_se), .CLK(CK), .Q(n3064), .QN(n1868) );
  SDFFX1 DFF_38_Q_reg ( .D(g8019), .SI(n3064), .SE(test_se), .CLK(CK), .Q(
        g4180), .QN() );
  SDFFX1 DFF_39_Q_reg ( .D(g6545), .SI(g4180), .SE(test_se), .CLK(CK), .Q(
        g1543), .QN() );
  SDFFX1 DFF_41_Q_reg ( .D(g256), .SI(g1543), .SE(test_se), .CLK(CK), .Q(g315), 
        .QN() );
  SDFFX1 DFF_42_Q_reg ( .D(g6533), .SI(g315), .SE(test_se), .CLK(CK), .Q(g1534), .QN(n1632) );
  SDFFX1 DFF_43_Q_reg ( .D(g8820), .SI(g1534), .SE(test_se), .CLK(CK), .Q(g622), .QN(n1713) );
  SDFFX1 DFF_44_Q_reg ( .D(g8941), .SI(g622), .SE(test_se), .CLK(CK), .Q(g1927), .QN() );
  SDFFX1 DFF_45_Q_reg ( .D(g10859), .SI(g1927), .SE(test_se), .CLK(CK), .Q(
        g1660), .QN() );
  SDFFX1 DFF_46_Q_reg ( .D(g6922), .SI(g1660), .SE(test_se), .CLK(CK), .Q(g278), .QN() );
  SDFFX1 DFF_47_Q_reg ( .D(g8772), .SI(g278), .SE(test_se), .CLK(CK), .Q(g1436), .QN() );
  SDFFX1 DFF_48_Q_reg ( .D(g8433), .SI(g1436), .SE(test_se), .CLK(CK), .Q(g718), .QN() );
  SDFFX1 DFF_49_Q_reg ( .D(g6526), .SI(g718), .SE(test_se), .CLK(CK), .Q(g8985), .QN(n1669) );
  SDFFX1 DFF_50_Q_reg ( .D(g10793), .SI(g8985), .SE(test_se), .CLK(CK), .Q(
        g554), .QN() );
  SDFFX1 DFF_51_Q_reg ( .D(g11333), .SI(g554), .SE(test_se), .CLK(CK), .Q(g496), .QN(n1689) );
  SDFFX1 DFF_52_Q_reg ( .D(g11392), .SI(g496), .SE(test_se), .CLK(CK), .Q(g981), .QN(n1720) );
  SDFFX1 DFF_53_Q_reg ( .D(n616), .SI(g981), .SE(test_se), .CLK(CK), .Q(g3007), 
        .QN(n1866) );
  SDFFX1 DFF_54_Q_reg ( .D(n1885), .SI(g3007), .SE(test_se), .CLK(CK), .Q(
        test_so1), .QN() );
  SDFFX1 DFF_55_Q_reg ( .D(g794), .SI(test_si2), .SE(test_se), .CLK(CK), .Q(
        g829), .QN(n1651) );
  SDFFX1 DFF_56_Q_reg ( .D(g6093), .SI(g829), .SE(test_se), .CLK(CK), .Q(g1095), .QN() );
  SDFFX1 DFF_57_Q_reg ( .D(g8889), .SI(g1095), .SE(test_se), .CLK(CK), .Q(g704), .QN() );
  SDFFX1 DFF_58_Q_reg ( .D(g7302), .SI(g704), .SE(test_se), .CLK(CK), .Q(g1265), .QN() );
  SDFFX1 DFF_59_Q_reg ( .D(g6525), .SI(g1265), .SE(test_se), .CLK(CK), .Q(
        g1786), .QN() );
  SDFFX1 DFF_60_Q_reg ( .D(g8429), .SI(g1786), .SE(test_se), .CLK(CK), .Q(g682), .QN() );
  SDFFX1 DFF_61_Q_reg ( .D(g7292), .SI(g682), .SE(test_se), .CLK(CK), .Q(g1296), .QN() );
  SDFFX1 DFF_62_Q_reg ( .D(g6284), .SI(g1296), .SE(test_se), .CLK(CK), .Q(
        g2602), .QN() );
  SDFFX1 DFF_63_Q_reg ( .D(g6621), .SI(g2602), .SE(test_se), .CLK(CK), .Q(
        g8977), .QN(n1668) );
  SDFFX1 DFF_64_Q_reg ( .D(g7134), .SI(g8977), .SE(test_se), .CLK(CK), .Q(
        n3062), .QN(n1595) );
  SDFFX1 DFF_65_Q_reg ( .D(g260), .SI(n3062), .SE(test_se), .CLK(CK), .Q(g327), 
        .QN() );
  SDFFX1 DFF_66_Q_reg ( .D(g6333), .SI(g327), .SE(test_se), .CLK(CK), .Q(g1389), .QN(n1603) );
  SDFFX1 DFF_67_Q_reg ( .D(g6826), .SI(g1389), .SE(test_se), .CLK(CK), .Q(
        g1371), .QN() );
  SDFFX1 DFF_68_Q_reg ( .D(g1955), .SI(g1371), .SE(test_se), .CLK(CK), .Q(
        g1956), .QN() );
  SDFFX1 DFF_69_Q_reg ( .D(g10860), .SI(g1956), .SE(test_se), .CLK(CK), .Q(
        g1675), .QN() );
  SDFFX1 DFF_70_Q_reg ( .D(g11483), .SI(g1675), .SE(test_se), .CLK(CK), .Q(
        g354), .QN() );
  SDFFX1 DFF_71_Q_reg ( .D(g6392), .SI(g354), .SE(test_se), .CLK(CK), .Q(g113), 
        .QN() );
  SDFFX1 DFF_72_Q_reg ( .D(g7626), .SI(g113), .SE(test_se), .CLK(CK), .Q(g639), 
        .QN(n1692) );
  SDFFX1 DFF_73_Q_reg ( .D(g10866), .SI(g639), .SE(test_se), .CLK(CK), .Q(
        g1684), .QN() );
  SDFFX1 DFF_74_Q_reg ( .D(g8193), .SI(g1684), .SE(test_se), .CLK(CK), .Q(
        g1639), .QN() );
  SDFFX1 DFF_75_Q_reg ( .D(g6983), .SI(g1639), .SE(test_se), .CLK(CK), .Q(
        g1791), .QN(n1702) );
  SDFFX1 DFF_76_Q_reg ( .D(g6839), .SI(g1791), .SE(test_se), .CLK(CK), .Q(g248), .QN(n1598) );
  SDFFX1 DFF_77_Q_reg ( .D(g4076), .SI(g248), .SE(test_se), .CLK(CK), .Q(g1707), .QN() );
  SDFFX1 DFF_78_Q_reg ( .D(g4293), .SI(g1707), .SE(test_se), .CLK(CK), .Q(
        g1759), .QN() );
  SDFFX1 DFF_79_Q_reg ( .D(g11482), .SI(g1759), .SE(test_se), .CLK(CK), .Q(
        g351), .QN() );
  SDFFX1 DFF_80_Q_reg ( .D(g1956), .SI(g351), .SE(test_se), .CLK(CK), .Q(g1957), .QN() );
  SDFFX1 DFF_81_Q_reg ( .D(g6507), .SI(g1957), .SE(test_se), .CLK(CK), .Q(
        g1604), .QN() );
  SDFFX1 DFF_82_Q_reg ( .D(g6096), .SI(g1604), .SE(test_se), .CLK(CK), .Q(
        g1098), .QN() );
  SDFFX1 DFF_83_Q_reg ( .D(g8250), .SI(g1098), .SE(test_se), .CLK(CK), .Q(g932), .QN(n1591) );
  SDFFX1 DFF_85_Q_reg ( .D(g8282), .SI(g932), .SE(test_se), .CLK(CK), .Q(g1896), .QN() );
  SDFFX1 DFF_86_Q_reg ( .D(g8435), .SI(g1896), .SE(test_se), .CLK(CK), .Q(g736), .QN() );
  SDFFX1 DFF_87_Q_reg ( .D(g6924), .SI(g736), .SE(test_se), .CLK(CK), .Q(g1019), .QN() );
  SDFFX1 DFF_88_Q_reg ( .D(g6819), .SI(g1019), .SE(test_se), .CLK(CK), .Q(
        n3061), .QN(n1625) );
  SDFFX1 DFF_89_Q_reg ( .D(g746), .SI(n3061), .SE(test_se), .CLK(CK), .Q(g745), 
        .QN() );
  SDFFX1 DFF_90_Q_reg ( .D(g6244), .SI(g745), .SE(test_se), .CLK(CK), .Q(g1419), .QN(n1602) );
  SDFFX1 DFF_91_Q_reg ( .D(g6627), .SI(g1419), .SE(test_se), .CLK(CK), .Q(
        g8979), .QN(n1667) );
  SDFFX1 DFF_92_Q_reg ( .D(n542), .SI(g8979), .SE(test_se), .CLK(CK), .Q(g32), 
        .QN() );
  SDFFX1 DFF_93_Q_reg ( .D(g3007), .SI(g32), .SE(test_se), .CLK(CK), .Q(n1865), 
        .QN() );
  SDFFX1 DFF_94_Q_reg ( .D(g6071), .SI(n1865), .SE(test_se), .CLK(CK), .Q(
        g1086), .QN() );
  SDFFX1 DFF_95_Q_reg ( .D(g8046), .SI(g1086), .SE(test_se), .CLK(CK), .Q(
        g1486), .QN() );
  SDFFX1 DFF_96_Q_reg ( .D(g10707), .SI(g1486), .SE(test_se), .CLK(CK), .Q(
        g1730), .QN() );
  SDFFX1 DFF_97_Q_reg ( .D(g6198), .SI(g1730), .SE(test_se), .CLK(CK), .Q(
        g1504), .QN() );
  SDFFX1 DFF_98_Q_reg ( .D(g8051), .SI(g1504), .SE(test_se), .CLK(CK), .Q(
        g1470), .QN() );
  SDFFX1 DFF_99_Q_reg ( .D(g8024), .SI(g1470), .SE(test_se), .CLK(CK), .Q(g822), .QN() );
  SDFFX1 DFF_100_Q_reg ( .D(g6253), .SI(g822), .SE(test_se), .CLK(CK), .Q(
        g2609), .QN() );
  SDFFX1 DFF_101_Q_reg ( .D(g10862), .SI(g2609), .SE(test_se), .CLK(CK), .Q(
        g1678), .QN() );
  SDFFX1 DFF_102_Q_reg ( .D(g8050), .SI(g1678), .SE(test_se), .CLK(CK), .Q(
        g174), .QN() );
  SDFFX1 DFF_103_Q_reg ( .D(g7133), .SI(g174), .SE(test_se), .CLK(CK), .Q(
        g1766), .QN() );
  SDFFX1 DFF_104_Q_reg ( .D(g7930), .SI(g1766), .SE(test_se), .CLK(CK), .Q(
        g1801), .QN() );
  SDFFX1 DFF_105_Q_reg ( .D(g6832), .SI(g1801), .SE(test_se), .CLK(CK), .Q(
        g186), .QN() );
  SDFFX1 DFF_106_Q_reg ( .D(g11308), .SI(g186), .SE(test_se), .CLK(CK), .Q(
        g959), .QN() );
  SDFFX1 DFF_108_Q_reg ( .D(g6918), .SI(g959), .SE(test_se), .CLK(CK), .Q(
        test_so2), .QN(n1869) );
  SDFFX1 DFF_109_Q_reg ( .D(g8769), .SI(test_si3), .SE(test_se), .CLK(CK), .Q(
        g1407), .QN() );
  SDFFX1 DFF_111_Q_reg ( .D(g6909), .SI(g1407), .SE(test_se), .CLK(CK), .Q(
        g1868), .QN() );
  SDFFX1 DFF_112_Q_reg ( .D(g4940), .SI(g1868), .SE(test_se), .CLK(CK), .Q(
        g4173), .QN() );
  SDFFX1 DFF_113_Q_reg ( .D(g5404), .SI(g4173), .SE(test_se), .CLK(CK), .Q(
        g1718), .QN(n1611) );
  SDFFX1 DFF_114_Q_reg ( .D(g11265), .SI(g1718), .SE(test_se), .CLK(CK), .Q(
        g396), .QN() );
  SDFFX1 DFF_115_Q_reg ( .D(g6930), .SI(g396), .SE(test_se), .CLK(CK), .Q(
        g1015), .QN() );
  SDFFX1 DFF_116_Q_reg ( .D(g10726), .SI(g1015), .SE(test_se), .CLK(CK), .Q(
        n1650), .QN() );
  SDFFX1 DFF_117_Q_reg ( .D(g4891), .SI(n1650), .SE(test_se), .CLK(CK), .Q(
        n3059), .QN(n1874) );
  SDFFX1 DFF_118_Q_reg ( .D(g6224), .SI(n3059), .SE(test_se), .CLK(CK), .Q(
        g1415), .QN() );
  SDFFX1 DFF_119_Q_reg ( .D(g7586), .SI(g1415), .SE(test_se), .CLK(CK), .Q(
        g1227), .QN() );
  SDFFX1 DFF_120_Q_reg ( .D(g10770), .SI(g1227), .SE(test_se), .CLK(CK), .Q(
        g1721), .QN() );
  SDFFX1 DFF_121_Q_reg ( .D(g2986), .SI(g1721), .SE(test_se), .CLK(CK), .Q(
        n3058), .QN(DFF_121_n1) );
  SDFFX1 DFF_122_Q_reg ( .D(n711), .SI(n3058), .SE(test_se), .CLK(CK), .Q(
        n3057), .QN(DFF_122_n1) );
  SDFFX1 DFF_123_Q_reg ( .D(g6934), .SI(n3057), .SE(test_se), .CLK(CK), .Q(
        g284), .QN() );
  SDFFX1 DFF_124_Q_reg ( .D(g11256), .SI(g284), .SE(test_se), .CLK(CK), .Q(
        g426), .QN() );
  SDFFX1 DFF_125_Q_reg ( .D(g6824), .SI(g426), .SE(test_se), .CLK(CK), .Q(g219), .QN() );
  SDFFX1 DFF_126_Q_reg ( .D(g1360), .SI(g219), .SE(test_se), .CLK(CK), .Q(
        n3056), .QN(DFF_126_n1) );
  SDFFX1 DFF_127_Q_reg ( .D(g6126), .SI(n3056), .SE(test_se), .CLK(CK), .Q(
        g806), .QN() );
  SDFFX1 DFF_128_Q_reg ( .D(g8767), .SI(g806), .SE(test_se), .CLK(CK), .Q(
        g1428), .QN() );
  SDFFX1 DFF_129_Q_reg ( .D(g6282), .SI(g1428), .SE(test_se), .CLK(CK), .Q(
        g2605), .QN() );
  SDFFX1 DFF_130_Q_reg ( .D(g6546), .SI(g2605), .SE(test_se), .CLK(CK), .Q(
        g1564), .QN() );
  SDFFX1 DFF_131_Q_reg ( .D(g4238), .SI(g1564), .SE(test_se), .CLK(CK), .Q(
        g1741), .QN(n1633) );
  SDFFX1 DFF_132_Q_reg ( .D(g6823), .SI(g1741), .SE(test_se), .CLK(CK), .Q(
        g225), .QN() );
  SDFFX1 DFF_133_Q_reg ( .D(g6928), .SI(g225), .SE(test_se), .CLK(CK), .Q(g281), .QN() );
  SDFFX1 DFF_134_Q_reg ( .D(g11602), .SI(g281), .SE(test_se), .CLK(CK), .Q(
        g1308), .QN() );
  SDFFX1 DFF_135_Q_reg ( .D(g9721), .SI(g1308), .SE(test_se), .CLK(CK), .Q(
        g611), .QN(n1609) );
  SDFFX1 DFF_136_Q_reg ( .D(g4890), .SI(g611), .SE(test_se), .CLK(CK), .Q(
        n3055), .QN(DFF_136_n1) );
  SDFFX1 DFF_137_Q_reg ( .D(n1586), .SI(n3055), .SE(test_se), .CLK(CK), .Q(
        g1217), .QN() );
  SDFFX1 DFF_138_Q_reg ( .D(g6524), .SI(g1217), .SE(test_se), .CLK(CK), .Q(
        g1589), .QN() );
  SDFFX1 DFF_139_Q_reg ( .D(g8045), .SI(g1589), .SE(test_se), .CLK(CK), .Q(
        g1466), .QN() );
  SDFFX1 DFF_140_Q_reg ( .D(g6469), .SI(g1466), .SE(test_se), .CLK(CK), .Q(
        g1571), .QN() );
  SDFFX1 DFF_141_Q_reg ( .D(g6471), .SI(g1571), .SE(test_se), .CLK(CK), .Q(
        g1861), .QN() );
  SDFFX1 DFF_142_Q_reg ( .D(g6821), .SI(g1861), .SE(test_se), .CLK(CK), .Q(
        n3054), .QN(n1688) );
  SDFFX1 DFF_143_Q_reg ( .D(g11514), .SI(n3054), .SE(test_se), .CLK(CK), .Q(
        g1448), .QN() );
  SDFFX1 DFF_145_Q_reg ( .D(g4480), .SI(g1448), .SE(test_se), .CLK(CK), .Q(
        g1133), .QN(n1706) );
  SDFFX1 DFF_146_Q_reg ( .D(g11610), .SI(g1133), .SE(test_se), .CLK(CK), .Q(
        g1333), .QN() );
  SDFFX1 DFF_147_Q_reg ( .D(g7843), .SI(g1333), .SE(test_se), .CLK(CK), .Q(
        g153), .QN() );
  SDFFX1 DFF_148_Q_reg ( .D(g11310), .SI(g153), .SE(test_se), .CLK(CK), .Q(
        g962), .QN(n1638) );
  SDFFX1 DFF_149_Q_reg ( .D(g5536), .SI(g962), .SE(test_se), .CLK(CK), .Q(
        g4175), .QN() );
  SDFFX1 DFF_150_Q_reg ( .D(g6285), .SI(g4175), .SE(test_se), .CLK(CK), .Q(
        g2603), .QN() );
  SDFFX1 DFF_151_Q_reg ( .D(g11331), .SI(g2603), .SE(test_se), .CLK(CK), .Q(
        g486), .QN(n1621) );
  SDFFX1 DFF_152_Q_reg ( .D(g11380), .SI(g486), .SE(test_se), .CLK(CK), .Q(
        g471), .QN(n1606) );
  SDFFX1 DFF_153_Q_reg ( .D(g6838), .SI(g471), .SE(test_se), .CLK(CK), .Q(
        g1397), .QN(n1711) );
  SDFFX1 DFF_154_Q_reg ( .D(g6283), .SI(g1397), .SE(test_se), .CLK(CK), .Q(
        g2606), .QN() );
  SDFFX1 DFF_155_Q_reg ( .D(g8288), .SI(g2606), .SE(test_se), .CLK(CK), .Q(
        g1950), .QN() );
  SDFFX1 DFF_156_Q_reg ( .D(g755), .SI(g1950), .SE(test_se), .CLK(CK), .Q(g756), .QN() );
  SDFFX1 DFF_157_Q_reg ( .D(g4892), .SI(g756), .SE(test_se), .CLK(CK), .Q(
        n3053), .QN(DFF_157_n1) );
  SDFFX1 DFF_159_Q_reg ( .D(g10855), .SI(g1101), .SE(test_se), .CLK(CK), .Q(
        g549), .QN() );
  SDFFX1 DFF_161_Q_reg ( .D(g10898), .SI(g549), .SE(test_se), .CLK(CK), .Q(
        g105), .QN() );
  SDFFX1 DFF_162_Q_reg ( .D(g10865), .SI(g105), .SE(test_se), .CLK(CK), .Q(
        g1669), .QN() );
  SDFFX1 DFF_163_Q_reg ( .D(g6822), .SI(g1669), .SE(test_se), .CLK(CK), .Q(
        test_so3), .QN() );
  SDFFX1 DFF_164_Q_reg ( .D(g6528), .SI(test_si4), .SE(test_se), .CLK(CK), .Q(
        g1531), .QN(n1652) );
  SDFFX1 DFF_165_Q_reg ( .D(g6180), .SI(g1531), .SE(test_se), .CLK(CK), .Q(
        g1458), .QN(n1703) );
  SDFFX1 DFF_166_Q_reg ( .D(g10718), .SI(g1458), .SE(test_se), .CLK(CK), .Q(
        g572), .QN() );
  SDFFX1 DFF_167_Q_reg ( .D(g6912), .SI(g572), .SE(test_se), .CLK(CK), .Q(
        g1011), .QN() );
  SDFFX1 DFF_168_Q_reg ( .D(g10719), .SI(g1011), .SE(test_se), .CLK(CK), .Q(
        n3051), .QN(DFF_168_n1) );
  SDFFX1 DFF_169_Q_reg ( .D(g6234), .SI(n3051), .SE(test_se), .CLK(CK), .Q(
        g1411), .QN() );
  SDFFX1 DFF_170_Q_reg ( .D(g6099), .SI(g1411), .SE(test_se), .CLK(CK), .Q(
        g1074), .QN() );
  SDFFX1 DFF_171_Q_reg ( .D(g11259), .SI(g1074), .SE(test_se), .CLK(CK), .Q(
        g444), .QN() );
  SDFFX1 DFF_172_Q_reg ( .D(g8039), .SI(g444), .SE(test_se), .CLK(CK), .Q(
        g1474), .QN() );
  SDFFX1 DFF_173_Q_reg ( .D(g6059), .SI(g1474), .SE(test_se), .CLK(CK), .Q(
        g1080), .QN() );
  SDFFX1 DFF_174_Q_reg ( .D(g5396), .SI(g1080), .SE(test_se), .CLK(CK), .Q(
        g1713), .QN(n1610) );
  SDFFX1 DFF_175_Q_reg ( .D(g262), .SI(g1713), .SE(test_se), .CLK(CK), .Q(g333), .QN() );
  SDFFX1 DFF_176_Q_reg ( .D(g6906), .SI(g333), .SE(test_se), .CLK(CK), .Q(g269), .QN() );
  SDFFX1 DFF_177_Q_reg ( .D(g11266), .SI(g269), .SE(test_se), .CLK(CK), .Q(
        g401), .QN() );
  SDFFX1 DFF_178_Q_reg ( .D(g11294), .SI(g401), .SE(test_se), .CLK(CK), .Q(
        g1857), .QN(n1682) );
  SDFFX1 DFF_179_Q_reg ( .D(g5421), .SI(g1857), .SE(test_se), .CLK(CK), .Q(g9), 
        .QN() );
  SDFFX1 DFF_180_Q_reg ( .D(g8649), .SI(g9), .SE(test_se), .CLK(CK), .Q(g664), 
        .QN() );
  SDFFX1 DFF_181_Q_reg ( .D(g11312), .SI(g664), .SE(test_se), .CLK(CK), .Q(
        g965), .QN(n1639) );
  SDFFX1 DFF_182_Q_reg ( .D(g6840), .SI(g965), .SE(test_se), .CLK(CK), .Q(
        g1400), .QN(n1629) );
  SDFFX1 DFF_183_Q_reg ( .D(g254), .SI(g1400), .SE(test_se), .CLK(CK), .Q(g309), .QN() );
  SDFFX1 DFF_184_Q_reg ( .D(g7202), .SI(g309), .SE(test_se), .CLK(CK), .Q(g814), .QN() );
  SDFFX1 DFF_185_Q_reg ( .D(g6834), .SI(g814), .SE(test_se), .CLK(CK), .Q(g231), .QN() );
  SDFFX1 DFF_186_Q_reg ( .D(g10795), .SI(g231), .SE(test_se), .CLK(CK), .Q(
        g557), .QN() );
  SDFFX1 DFF_187_Q_reg ( .D(g6283), .SI(g557), .SE(test_se), .CLK(CK), .Q(
        g2612), .QN() );
  SDFFX1 DFF_188_Q_reg ( .D(g875), .SI(g2612), .SE(test_se), .CLK(CK), .Q(g869), .QN() );
  SDFFX1 DFF_189_Q_reg ( .D(g6831), .SI(g869), .SE(test_se), .CLK(CK), .Q(
        g1383), .QN() );
  SDFFX1 DFF_190_Q_reg ( .D(g8060), .SI(g1383), .SE(test_se), .CLK(CK), .Q(
        g158), .QN() );
  SDFFX1 DFF_191_Q_reg ( .D(g4893), .SI(g158), .SE(test_se), .CLK(CK), .Q(g627), .QN(n1701) );
  SDFFX1 DFF_192_Q_reg ( .D(g7244), .SI(g627), .SE(test_se), .CLK(CK), .Q(
        g1023), .QN() );
  SDFFX1 DFF_193_Q_reg ( .D(g6026), .SI(g1023), .SE(test_se), .CLK(CK), .Q(
        g259), .QN() );
  SDFFX1 DFF_194_Q_reg ( .D(g3069), .SI(g259), .SE(test_se), .CLK(CK), .Q(
        n3050), .QN(DFF_194_n1) );
  SDFFX1 DFF_195_Q_reg ( .D(g11608), .SI(n3050), .SE(test_se), .CLK(CK), .Q(
        g1327), .QN() );
  SDFFX1 DFF_196_Q_reg ( .D(g7660), .SI(g1327), .SE(test_se), .CLK(CK), .Q(
        g654), .QN() );
  SDFFX1 DFF_197_Q_reg ( .D(g6911), .SI(g654), .SE(test_se), .CLK(CK), .Q(g293), .QN() );
  SDFFX1 DFF_198_Q_reg ( .D(g11640), .SI(g293), .SE(test_se), .CLK(CK), .Q(
        g1346), .QN() );
  SDFFX1 DFF_199_Q_reg ( .D(g8777), .SI(g1346), .SE(test_se), .CLK(CK), .Q(
        g1633), .QN() );
  SDFFX1 DFF_200_Q_reg ( .D(g4274), .SI(g1633), .SE(test_se), .CLK(CK), .Q(
        g1753), .QN() );
  SDFFX1 DFF_201_Q_reg ( .D(n518), .SI(g1753), .SE(test_se), .CLK(CK), .Q(
        g1508), .QN(n1707) );
  SDFFX1 DFF_202_Q_reg ( .D(g7297), .SI(g1508), .SE(test_se), .CLK(CK), .Q(
        g1240), .QN() );
  SDFFX1 DFF_203_Q_reg ( .D(g11326), .SI(g1240), .SE(test_se), .CLK(CK), .Q(
        g538), .QN() );
  SDFFX1 DFF_204_Q_reg ( .D(g11269), .SI(g538), .SE(test_se), .CLK(CK), .Q(
        g416), .QN() );
  SDFFX1 DFF_205_Q_reg ( .D(g11325), .SI(g416), .SE(test_se), .CLK(CK), .Q(
        g542), .QN() );
  SDFFX1 DFF_206_Q_reg ( .D(g10864), .SI(g542), .SE(test_se), .CLK(CK), .Q(
        g1681), .QN() );
  SDFFX1 DFF_207_Q_reg ( .D(g11290), .SI(g1681), .SE(test_se), .CLK(CK), .Q(
        g374), .QN() );
  SDFFX1 DFF_208_Q_reg ( .D(g10798), .SI(g374), .SE(test_se), .CLK(CK), .Q(
        g563), .QN() );
  SDFFX1 DFF_209_Q_reg ( .D(g8284), .SI(g563), .SE(test_se), .CLK(CK), .Q(
        g1914), .QN() );
  SDFFX1 DFF_210_Q_reg ( .D(g11328), .SI(g1914), .SE(test_se), .CLK(CK), .Q(
        g530), .QN() );
  SDFFX1 DFF_211_Q_reg ( .D(g10800), .SI(g530), .SE(test_se), .CLK(CK), .Q(
        g575), .QN() );
  SDFFX1 DFF_212_Q_reg ( .D(g8944), .SI(g575), .SE(test_se), .CLK(CK), .Q(
        g1936), .QN(n1694) );
  SDFFX1 DFF_213_Q_reg ( .D(g7183), .SI(g1936), .SE(test_se), .CLK(CK), .Q(
        g8978), .QN(n1674) );
  SDFFX1 DFF_214_Q_reg ( .D(g4465), .SI(g8978), .SE(test_se), .CLK(CK), .Q(
        test_so4), .QN(n1661) );
  SDFFX1 DFF_215_Q_reg ( .D(g1356), .SI(test_si5), .SE(test_se), .CLK(CK), .Q(
        g1317), .QN() );
  SDFFX1 DFF_216_Q_reg ( .D(g11484), .SI(g1317), .SE(test_se), .CLK(CK), .Q(
        g357), .QN() );
  SDFFX1 DFF_217_Q_reg ( .D(g11263), .SI(g357), .SE(test_se), .CLK(CK), .Q(
        g386), .QN() );
  SDFFX1 DFF_218_Q_reg ( .D(g6501), .SI(g386), .SE(test_se), .CLK(CK), .Q(
        g1601), .QN() );
  SDFFX1 DFF_220_Q_reg ( .D(g6757), .SI(g1601), .SE(test_se), .CLK(CK), .Q(
        g166), .QN() );
  SDFFX1 DFF_221_Q_reg ( .D(g11334), .SI(g166), .SE(test_se), .CLK(CK), .Q(
        g501), .QN(n1690) );
  SDFFX1 DFF_222_Q_reg ( .D(g6042), .SI(g501), .SE(test_se), .CLK(CK), .Q(g262), .QN() );
  SDFFX1 DFF_223_Q_reg ( .D(g8384), .SI(g262), .SE(test_se), .CLK(CK), .Q(
        g1840), .QN() );
  SDFFX1 DFF_224_Q_reg ( .D(g6653), .SI(g1840), .SE(test_se), .CLK(CK), .Q(
        g8983), .QN(n1666) );
  SDFFX1 DFF_225_Q_reg ( .D(g257), .SI(g8983), .SE(test_se), .CLK(CK), .Q(g318), .QN() );
  SDFFX1 DFF_226_Q_reg ( .D(g5763), .SI(g318), .SE(test_se), .CLK(CK), .Q(
        g1356), .QN() );
  SDFFX1 DFF_227_Q_reg ( .D(g5849), .SI(g1356), .SE(test_se), .CLK(CK), .Q(
        g794), .QN() );
  SDFFX1 DFF_228_Q_reg ( .D(g10722), .SI(g794), .SE(test_se), .CLK(CK), .Q(
        n3048), .QN(DFF_228_n1) );
  SDFFX1 DFF_229_Q_reg ( .D(g6929), .SI(n3048), .SE(test_se), .CLK(CK), .Q(
        g302), .QN() );
  SDFFX1 DFF_230_Q_reg ( .D(g11488), .SI(g302), .SE(test_se), .CLK(CK), .Q(
        g342), .QN() );
  SDFFX1 DFF_231_Q_reg ( .D(g7299), .SI(g342), .SE(test_se), .CLK(CK), .Q(
        g1250), .QN() );
  SDFFX1 DFF_232_Q_reg ( .D(g4330), .SI(g1250), .SE(test_se), .CLK(CK), .Q(
        g1163), .QN() );
  SDFFX1 DFF_233_Q_reg ( .D(g1958), .SI(g1163), .SE(test_se), .CLK(CK), .Q(
        n3047), .QN(g8271) );
  SDFFX1 DFF_234_Q_reg ( .D(g7257), .SI(n3047), .SE(test_se), .CLK(CK), .Q(
        g1032), .QN() );
  SDFFX1 DFF_235_Q_reg ( .D(g8775), .SI(g1032), .SE(test_se), .CLK(CK), .Q(
        g1432), .QN() );
  SDFFX1 DFF_237_Q_reg ( .D(g5770), .SI(g1432), .SE(test_se), .CLK(CK), .Q(
        g1453), .QN(n1628) );
  SDFFX1 DFF_238_Q_reg ( .D(g11486), .SI(g1453), .SE(test_se), .CLK(CK), .Q(
        g363), .QN() );
  SDFFX1 DFF_239_Q_reg ( .D(g261), .SI(g363), .SE(test_se), .CLK(CK), .Q(g330), 
        .QN() );
  SDFFX1 DFF_240_Q_reg ( .D(g4338), .SI(g330), .SE(test_se), .CLK(CK), .Q(
        g1157), .QN() );
  SDFFX1 DFF_241_Q_reg ( .D(g4500), .SI(g1157), .SE(test_se), .CLK(CK), .Q(
        n3046), .QN(n1648) );
  SDFFX1 DFF_242_Q_reg ( .D(g10721), .SI(n3046), .SE(test_se), .CLK(CK), .Q(
        n3045), .QN(DFF_242_n1) );
  SDFFX1 DFF_243_Q_reg ( .D(g8147), .SI(n3045), .SE(test_se), .CLK(CK), .Q(
        g928), .QN(n1604) );
  SDFFX1 DFF_244_Q_reg ( .D(g6038), .SI(g928), .SE(test_se), .CLK(CK), .Q(g261), .QN() );
  SDFFX1 DFF_245_Q_reg ( .D(g11337), .SI(g261), .SE(test_se), .CLK(CK), .Q(
        g516), .QN(n1620) );
  SDFFX1 DFF_246_Q_reg ( .D(g6045), .SI(g516), .SE(test_se), .CLK(CK), .Q(g254), .QN() );
  SDFFX1 DFF_247_Q_reg ( .D(g7191), .SI(g254), .SE(test_se), .CLK(CK), .Q(
        g4178), .QN() );
  SDFFX1 DFF_248_Q_reg ( .D(g826), .SI(g4178), .SE(test_se), .CLK(CK), .Q(g861), .QN() );
  SDFFX1 DFF_249_Q_reg ( .D(g8774), .SI(g861), .SE(test_se), .CLK(CK), .Q(
        g1627), .QN() );
  SDFFX1 DFF_250_Q_reg ( .D(g7293), .SI(g1627), .SE(test_se), .CLK(CK), .Q(
        g1292), .QN() );
  SDFFX1 DFF_251_Q_reg ( .D(g6907), .SI(g1292), .SE(test_se), .CLK(CK), .Q(
        g290), .QN() );
  SDFFX1 DFF_252_Q_reg ( .D(g4903), .SI(g290), .SE(test_se), .CLK(CK), .Q(
        n3044), .QN(n1873) );
  SDFFX1 DFF_253_Q_reg ( .D(g6123), .SI(n3044), .SE(test_se), .CLK(CK), .Q(
        g4176), .QN() );
  SDFFX1 DFF_254_Q_reg ( .D(g6506), .SI(g4176), .SE(test_se), .CLK(CK), .Q(
        g1583), .QN() );
  SDFFX1 DFF_255_Q_reg ( .D(g11376), .SI(g1583), .SE(test_se), .CLK(CK), .Q(
        g466), .QN(n1646) );
  SDFFX1 DFF_256_Q_reg ( .D(g6542), .SI(g466), .SE(test_se), .CLK(CK), .Q(
        g1561), .QN() );
  SDFFX1 DFF_258_Q_reg ( .D(g6551), .SI(g1561), .SE(test_se), .CLK(CK), .Q(
        g1546), .QN() );
  SDFFX1 DFF_259_Q_reg ( .D(g6901), .SI(g1546), .SE(test_se), .CLK(CK), .Q(
        g287), .QN() );
  SDFFX1 DFF_260_Q_reg ( .D(g10797), .SI(g287), .SE(test_se), .CLK(CK), .Q(
        g560), .QN() );
  SDFFX1 DFF_261_Q_reg ( .D(g8505), .SI(g560), .SE(test_se), .CLK(CK), .Q(g617), .QN(n1645) );
  SDFFX1 DFF_262_Q_reg ( .D(n667), .SI(g617), .SE(test_se), .CLK(CK), .Q(n1631), .QN() );
  SDFFX1 DFF_263_Q_reg ( .D(g11647), .SI(n1631), .SE(test_se), .CLK(CK), .Q(
        g336), .QN() );
  SDFFX1 DFF_264_Q_reg ( .D(g11340), .SI(g336), .SE(test_se), .CLK(CK), .Q(
        g456), .QN(n1641) );
  SDFFX1 DFF_265_Q_reg ( .D(g253), .SI(g456), .SE(test_se), .CLK(CK), .Q(g305), 
        .QN(n1681) );
  SDFFX1 DFF_266_Q_reg ( .D(g11625), .SI(g305), .SE(test_se), .CLK(CK), .Q(
        g345), .QN() );
  SDFFX1 DFF_267_Q_reg ( .D(g636), .SI(g345), .SE(test_se), .CLK(CK), .Q(g8), 
        .QN() );
  SDFFX1 DFF_268_Q_reg ( .D(g6502), .SI(g8), .SE(test_se), .CLK(CK), .Q(
        test_so5), .QN() );
  SDFFX1 DFF_269_Q_reg ( .D(N599), .SI(test_si6), .SE(test_se), .CLK(CK), .Q(
        g2648), .QN() );
  SDFFX1 DFF_270_Q_reg ( .D(g6049), .SI(g2648), .SE(test_se), .CLK(CK), .Q(
        g255), .QN() );
  SDFFX1 DFF_271_Q_reg ( .D(g8945), .SI(g255), .SE(test_se), .CLK(CK), .Q(
        g1945), .QN(n1697) );
  SDFFX1 DFF_272_Q_reg ( .D(g4231), .SI(g1945), .SE(test_se), .CLK(CK), .Q(
        g1738), .QN(n1640) );
  SDFFX1 DFF_273_Q_reg ( .D(g8040), .SI(g1738), .SE(test_se), .CLK(CK), .Q(
        g1478), .QN() );
  SDFFX1 DFF_275_Q_reg ( .D(n562), .SI(g1478), .SE(test_se), .CLK(CK), .Q(
        n3042), .QN(DFF_275_n1) );
  SDFFX1 DFF_276_Q_reg ( .D(g6155), .SI(n3042), .SE(test_se), .CLK(CK), .Q(
        g1690), .QN(n1653) );
  SDFFX1 DFF_277_Q_reg ( .D(g8043), .SI(g1690), .SE(test_se), .CLK(CK), .Q(
        g1482), .QN() );
  SDFFX1 DFF_278_Q_reg ( .D(g5173), .SI(g1482), .SE(test_se), .CLK(CK), .Q(
        g1110), .QN(n1677) );
  SDFFX1 DFF_279_Q_reg ( .D(g6916), .SI(g1110), .SE(test_se), .CLK(CK), .Q(
        g296), .QN() );
  SDFFX1 DFF_280_Q_reg ( .D(g10861), .SI(g296), .SE(test_se), .CLK(CK), .Q(
        g1663), .QN() );
  SDFFX1 DFF_281_Q_reg ( .D(g8431), .SI(g1663), .SE(test_se), .CLK(CK), .Q(
        g700), .QN() );
  SDFFX1 DFF_282_Q_reg ( .D(g4309), .SI(g700), .SE(test_se), .CLK(CK), .Q(
        g1762), .QN() );
  SDFFX1 DFF_283_Q_reg ( .D(g11485), .SI(g1762), .SE(test_se), .CLK(CK), .Q(
        g360), .QN() );
  SDFFX1 DFF_284_Q_reg ( .D(g6334), .SI(g360), .SE(test_se), .CLK(CK), .Q(g192), .QN() );
  SDFFX1 DFF_285_Q_reg ( .D(g10767), .SI(g192), .SE(test_se), .CLK(CK), .Q(
        g1657), .QN() );
  SDFFX1 DFF_286_Q_reg ( .D(g8923), .SI(g1657), .SE(test_se), .CLK(CK), .Q(
        g722), .QN(n1693) );
  SDFFX1 DFF_287_Q_reg ( .D(g7189), .SI(g722), .SE(test_se), .CLK(CK), .Q(
        g8980), .QN(n1673) );
  SDFFX1 DFF_288_Q_reg ( .D(g10799), .SI(g8980), .SE(test_se), .CLK(CK), .Q(
        g566), .QN() );
  SDFFX1 DFF_289_Q_reg ( .D(g6747), .SI(g566), .SE(test_se), .CLK(CK), .Q(
        n3041), .QN(n1714) );
  SDFFX1 DFF_290_Q_reg ( .D(g6080), .SI(n3041), .SE(test_se), .CLK(CK), .Q(
        g1089), .QN() );
  SDFFX1 DFF_291_Q_reg ( .D(g3381), .SI(g1089), .SE(test_se), .CLK(CK), .Q(
        g2986), .QN() );
  SDFFX1 DFF_292_Q_reg ( .D(g5910), .SI(g2986), .SE(test_se), .CLK(CK), .Q(
        g1071), .QN() );
  SDFFX1 DFF_293_Q_reg ( .D(g11393), .SI(g1071), .SE(test_se), .CLK(CK), .Q(
        g986), .QN(n1722) );
  SDFFX1 DFF_294_Q_reg ( .D(g11349), .SI(g986), .SE(test_se), .CLK(CK), .Q(
        g971), .QN() );
  SDFFX1 DFF_295_Q_reg ( .D(g6265), .SI(g971), .SE(test_se), .CLK(CK), .Q(
        g1955), .QN() );
  SDFFX1 DFF_296_Q_reg ( .D(g6439), .SI(g1955), .SE(test_se), .CLK(CK), .Q(
        g143), .QN() );
  SDFFX1 DFF_297_Q_reg ( .D(g9266), .SI(g143), .SE(test_se), .CLK(CK), .Q(
        g1814), .QN(n1608) );
  SDFFX1 DFF_299_Q_reg ( .D(g1217), .SI(g1814), .SE(test_se), .CLK(CK), .Q(
        g1212), .QN() );
  SDFFX1 DFF_300_Q_reg ( .D(g8940), .SI(g1212), .SE(test_se), .CLK(CK), .Q(
        g1918), .QN() );
  SDFFX1 DFF_301_Q_reg ( .D(g7705), .SI(g1918), .SE(test_se), .CLK(CK), .Q(
        g4179), .QN() );
  SDFFX1 DFF_302_Q_reg ( .D(g9269), .SI(g4179), .SE(test_se), .CLK(CK), .Q(
        g1822), .QN(n1643) );
  SDFFX1 DFF_303_Q_reg ( .D(g6820), .SI(g1822), .SE(test_se), .CLK(CK), .Q(
        g237), .QN() );
  SDFFX1 DFF_304_Q_reg ( .D(g756), .SI(g237), .SE(test_se), .CLK(CK), .Q(g746), 
        .QN() );
  SDFFX1 DFF_306_Q_reg ( .D(g8042), .SI(g746), .SE(test_se), .CLK(CK), .Q(
        g1462), .QN() );
  SDFFX1 DFF_307_Q_reg ( .D(g6759), .SI(g1462), .SE(test_se), .CLK(CK), .Q(
        g178), .QN() );
  SDFFX1 DFF_308_Q_reg ( .D(g11487), .SI(g178), .SE(test_se), .CLK(CK), .Q(
        g366), .QN() );
  SDFFX1 DFF_309_Q_reg ( .D(g802), .SI(g366), .SE(test_se), .CLK(CK), .Q(g837), 
        .QN() );
  SDFFX1 DFF_310_Q_reg ( .D(g9124), .SI(g837), .SE(test_se), .CLK(CK), .Q(g599), .QN(n1644) );
  SDFFX1 DFF_311_Q_reg ( .D(g11293), .SI(g599), .SE(test_se), .CLK(CK), .Q(
        g1854), .QN(DFF_311_n1) );
  SDFFX1 DFF_312_Q_reg ( .D(g11298), .SI(g1854), .SE(test_se), .CLK(CK), .Q(
        g944), .QN() );
  SDFFX1 DFF_313_Q_reg ( .D(g8287), .SI(g944), .SE(test_se), .CLK(CK), .Q(
        g1941), .QN() );
  SDFFX1 DFF_314_Q_reg ( .D(g8047), .SI(g1941), .SE(test_se), .CLK(CK), .Q(
        g170), .QN() );
  SDFFX1 DFF_315_Q_reg ( .D(g6205), .SI(g170), .SE(test_se), .CLK(CK), .Q(
        g1520), .QN(n1710) );
  SDFFX1 DFF_316_Q_reg ( .D(g8885), .SI(g1520), .SE(test_se), .CLK(CK), .Q(
        g686), .QN(n1676) );
  SDFFX1 DFF_317_Q_reg ( .D(g11305), .SI(g686), .SE(test_se), .CLK(CK), .Q(
        g953), .QN() );
  SDFFX1 DFF_318_Q_reg ( .D(g5556), .SI(g953), .SE(test_se), .CLK(CK), .Q(
        g1958), .QN() );
  SDFFX1 DFF_319_Q_reg ( .D(g10664), .SI(g1958), .SE(test_se), .CLK(CK), .Q(
        n3040), .QN(DFF_319_n1) );
  SDFFX1 DFF_320_Q_reg ( .D(g2478), .SI(n3040), .SE(test_se), .CLK(CK), .Q(
        g1765), .QN() );
  SDFFX1 DFF_321_Q_reg ( .D(g10711), .SI(g1765), .SE(test_se), .CLK(CK), .Q(
        g1733), .QN() );
  SDFFX1 DFF_322_Q_reg ( .D(g7303), .SI(g1733), .SE(test_se), .CLK(CK), .Q(
        test_so6), .QN() );
  SDFFX1 DFF_323_Q_reg ( .D(g5194), .SI(test_si7), .SE(test_se), .CLK(CK), .Q(
        g1610), .QN() );
  SDFFX1 DFF_324_Q_reg ( .D(g7541), .SI(g1610), .SE(test_se), .CLK(CK), .Q(
        g1796), .QN(n1626) );
  SDFFX1 DFF_325_Q_reg ( .D(g11607), .SI(g1796), .SE(test_se), .CLK(CK), .Q(
        g1324), .QN() );
  SDFFX1 DFF_326_Q_reg ( .D(g6541), .SI(g1324), .SE(test_se), .CLK(CK), .Q(
        g1540), .QN() );
  SDFFX1 DFF_327_Q_reg ( .D(g6827), .SI(g1540), .SE(test_se), .CLK(CK), .Q(
        n3038), .QN(n1624) );
  SDFFX1 DFF_328_Q_reg ( .D(n687), .SI(n3038), .SE(test_se), .CLK(CK), .Q(
        g3069), .QN() );
  SDFFX1 DFF_329_Q_reg ( .D(g11332), .SI(g3069), .SE(test_se), .CLK(CK), .Q(
        g491), .QN(n1691) );
  SDFFX1 DFF_330_Q_reg ( .D(g4902), .SI(g491), .SE(test_se), .CLK(CK), .Q(
        n3037), .QN(DFF_330_n1) );
  SDFFX1 DFF_331_Q_reg ( .D(g6828), .SI(n3037), .SE(test_se), .CLK(CK), .Q(
        g213), .QN() );
  SDFFX1 DFF_332_Q_reg ( .D(g6516), .SI(g213), .SE(test_se), .CLK(CK), .Q(
        g1781), .QN(n1659) );
  SDFFX1 DFF_333_Q_reg ( .D(g8938), .SI(g1781), .SE(test_se), .CLK(CK), .Q(
        g1900), .QN(n1675) );
  SDFFX1 DFF_334_Q_reg ( .D(g7298), .SI(g1900), .SE(test_se), .CLK(CK), .Q(
        g1245), .QN() );
  SDFFX1 DFF_335_Q_reg ( .D(n550), .SI(g1245), .SE(test_se), .CLK(CK), .Q(
        n3036), .QN(n1683) );
  SDFFX1 DFF_336_Q_reg ( .D(g6672), .SI(n3036), .SE(test_se), .CLK(CK), .Q(
        n3035), .QN(DFF_336_n1) );
  SDFFX1 DFF_337_Q_reg ( .D(g8048), .SI(n3035), .SE(test_se), .CLK(CK), .Q(
        g148), .QN() );
  SDFFX1 DFF_338_Q_reg ( .D(g798), .SI(g148), .SE(test_se), .CLK(CK), .Q(g833), 
        .QN() );
  SDFFX1 DFF_339_Q_reg ( .D(g8285), .SI(g833), .SE(test_se), .CLK(CK), .Q(
        g1923), .QN(n1718) );
  SDFFX1 DFF_340_Q_reg ( .D(g8254), .SI(g1923), .SE(test_se), .CLK(CK), .Q(
        g936), .QN(n1630) );
  SDFFX1 DFF_342_Q_reg ( .D(g11604), .SI(g936), .SE(test_se), .CLK(CK), .Q(
        g1314), .QN() );
  SDFFX1 DFF_343_Q_reg ( .D(g814), .SI(g1314), .SE(test_se), .CLK(CK), .Q(g849), .QN() );
  SDFFX1 DFF_344_Q_reg ( .D(g11636), .SI(g849), .SE(test_se), .CLK(CK), .Q(
        g1336), .QN() );
  SDFFX1 DFF_345_Q_reg ( .D(g6910), .SI(g1336), .SE(test_se), .CLK(CK), .Q(
        g272), .QN() );
  SDFFX1 DFF_346_Q_reg ( .D(g8173), .SI(g272), .SE(test_se), .CLK(CK), .Q(
        g1806), .QN() );
  SDFFX1 DFF_347_Q_reg ( .D(g8245), .SI(g1806), .SE(test_se), .CLK(CK), .Q(
        g826), .QN(n1716) );
  SDFFX1 DFF_349_Q_reg ( .D(g8281), .SI(g826), .SE(test_se), .CLK(CK), .Q(
        g1887), .QN() );
  SDFFX1 DFF_350_Q_reg ( .D(g10724), .SI(g1887), .SE(test_se), .CLK(CK), .Q(
        n3034), .QN(DFF_350_n1) );
  SDFFX1 DFF_351_Q_reg ( .D(g11314), .SI(n3034), .SE(test_se), .CLK(CK), .Q(
        g968), .QN() );
  SDFFX1 DFF_352_Q_reg ( .D(g4905), .SI(g968), .SE(test_se), .CLK(CK), .Q(
        n3033), .QN(n1642) );
  SDFFX1 DFF_353_Q_reg ( .D(g4484), .SI(n3033), .SE(test_se), .CLK(CK), .Q(
        g1137), .QN(n1597) );
  SDFFX1 DFF_354_Q_reg ( .D(g8937), .SI(g1137), .SE(test_se), .CLK(CK), .Q(
        g1891), .QN(n1657) );
  SDFFX1 DFF_355_Q_reg ( .D(g7300), .SI(g1891), .SE(test_se), .CLK(CK), .Q(
        g1255), .QN() );
  SDFFX1 DFF_356_Q_reg ( .D(g6002), .SI(g1255), .SE(test_se), .CLK(CK), .Q(
        g257), .QN() );
  SDFFX1 DFF_357_Q_reg ( .D(n1588), .SI(g257), .SE(test_se), .CLK(CK), .Q(g874), .QN() );
  SDFFX1 DFF_358_Q_reg ( .D(g9110), .SI(g874), .SE(test_se), .CLK(CK), .Q(g591), .QN(n1607) );
  SDFFX1 DFF_359_Q_reg ( .D(g8926), .SI(g591), .SE(test_se), .CLK(CK), .Q(g731), .QN(n1696) );
  SDFFX1 DFF_360_Q_reg ( .D(g8631), .SI(g731), .SE(test_se), .CLK(CK), .Q(g636), .QN() );
  SDFFX1 DFF_361_Q_reg ( .D(g7632), .SI(g636), .SE(test_se), .CLK(CK), .Q(
        g1218), .QN() );
  SDFFX1 DFF_362_Q_reg ( .D(g9150), .SI(g1218), .SE(test_se), .CLK(CK), .Q(
        g605), .QN(n1593) );
  SDFFX1 DFF_363_Q_reg ( .D(g6531), .SI(g605), .SE(test_se), .CLK(CK), .Q(
        g8986), .QN(n1665) );
  SDFFX1 DFF_364_Q_reg ( .D(g6786), .SI(g8986), .SE(test_se), .CLK(CK), .Q(
        g182), .QN() );
  SDFFX1 DFF_365_Q_reg ( .D(g11303), .SI(g182), .SE(test_se), .CLK(CK), .Q(
        g950), .QN() );
  SDFFX1 DFF_366_Q_reg ( .D(g4477), .SI(g950), .SE(test_se), .CLK(CK), .Q(
        g1129), .QN(n1705) );
  SDFFX1 DFF_367_Q_reg ( .D(g822), .SI(g1129), .SE(test_se), .CLK(CK), .Q(g857), .QN() );
  SDFFX1 DFF_368_Q_reg ( .D(g11258), .SI(g857), .SE(test_se), .CLK(CK), .Q(
        g448), .QN() );
  SDFFX1 DFF_369_Q_reg ( .D(g9272), .SI(g448), .SE(test_se), .CLK(CK), .Q(
        g1828), .QN(n1605) );
  SDFFX1 DFF_370_Q_reg ( .D(g10773), .SI(g1828), .SE(test_se), .CLK(CK), .Q(
        g1727), .QN() );
  SDFFX1 DFF_371_Q_reg ( .D(g6470), .SI(g1727), .SE(test_se), .CLK(CK), .Q(
        g1592), .QN() );
  SDFFX1 DFF_372_Q_reg ( .D(g5083), .SI(g1592), .SE(test_se), .CLK(CK), .Q(
        g1703), .QN() );
  SDFFX1 DFF_373_Q_reg ( .D(g8286), .SI(g1703), .SE(test_se), .CLK(CK), .Q(
        g1932), .QN() );
  SDFFX1 DFF_374_Q_reg ( .D(g8773), .SI(g1932), .SE(test_se), .CLK(CK), .Q(
        g1624), .QN() );
  SDFFX1 DFF_376_Q_reg ( .D(g6054), .SI(g1624), .SE(test_se), .CLK(CK), .Q(
        test_so7), .QN() );
  SDFFX1 DFF_377_Q_reg ( .D(g6281), .SI(test_si8), .SE(test_se), .CLK(CK), .Q(
        g2601), .QN() );
  SDFFX1 DFF_378_Q_reg ( .D(g11260), .SI(g2601), .SE(test_se), .CLK(CK), .Q(
        g440), .QN() );
  SDFFX1 DFF_379_Q_reg ( .D(g11338), .SI(g440), .SE(test_se), .CLK(CK), .Q(
        g476), .QN(n1599) );
  SDFFX1 DFF_380_Q_reg ( .D(g5918), .SI(g476), .SE(test_se), .CLK(CK), .Q(g119), .QN(n1613) );
  SDFFX1 DFF_381_Q_reg ( .D(g8922), .SI(g119), .SE(test_se), .CLK(CK), .Q(g668), .QN(n1662) );
  SDFFX1 DFF_382_Q_reg ( .D(g8049), .SI(g668), .SE(test_se), .CLK(CK), .Q(g139), .QN() );
  SDFFX1 DFF_383_Q_reg ( .D(g4342), .SI(g139), .SE(test_se), .CLK(CK), .Q(
        g1149), .QN(n1685) );
  SDFFX1 DFF_384_Q_reg ( .D(g10720), .SI(g1149), .SE(test_se), .CLK(CK), .Q(
        n3031), .QN(DFF_384_n1) );
  SDFFX1 DFF_385_Q_reg ( .D(g6755), .SI(n3031), .SE(test_se), .CLK(CK), .Q(
        n3030), .QN(DFF_385_n1) );
  SDFFX1 DFF_386_Q_reg ( .D(g6897), .SI(n3030), .SE(test_se), .CLK(CK), .Q(
        g263), .QN() );
  SDFFX1 DFF_387_Q_reg ( .D(g7709), .SI(g263), .SE(test_se), .CLK(CK), .Q(g818), .QN() );
  SDFFX1 DFF_388_Q_reg ( .D(g4255), .SI(g818), .SE(test_se), .CLK(CK), .Q(
        g1747), .QN() );
  SDFFX1 DFF_389_Q_reg ( .D(g5543), .SI(g1747), .SE(test_se), .CLK(CK), .Q(
        g802), .QN(n1622) );
  SDFFX1 DFF_390_Q_reg ( .D(g6915), .SI(g802), .SE(test_se), .CLK(CK), .Q(g275), .QN() );
  SDFFX1 DFF_391_Q_reg ( .D(g6513), .SI(g275), .SE(test_se), .CLK(CK), .Q(
        g1524), .QN(n1649) );
  SDFFX1 DFF_392_Q_reg ( .D(g6480), .SI(g1524), .SE(test_se), .CLK(CK), .Q(
        g1577), .QN() );
  SDFFX1 DFF_393_Q_reg ( .D(g6733), .SI(g1577), .SE(test_se), .CLK(CK), .Q(
        g810), .QN() );
  SDFFX1 DFF_394_Q_reg ( .D(g11264), .SI(g810), .SE(test_se), .CLK(CK), .Q(
        g391), .QN() );
  SDFFX1 DFF_395_Q_reg ( .D(g8973), .SI(g391), .SE(test_se), .CLK(CK), .Q(g658), .QN(n1615) );
  SDFFX1 DFF_396_Q_reg ( .D(g6833), .SI(g658), .SE(test_se), .CLK(CK), .Q(
        g1386), .QN() );
  SDFFX1 DFF_397_Q_reg ( .D(g5996), .SI(g1386), .SE(test_se), .CLK(CK), .Q(
        g253), .QN() );
  SDFFX1 DFF_398_Q_reg ( .D(n1587), .SI(g253), .SE(test_se), .CLK(CK), .Q(g875), .QN() );
  SDFFX1 DFF_399_Q_reg ( .D(g4473), .SI(g875), .SE(test_se), .CLK(CK), .Q(
        g1125), .QN(n1708) );
  SDFFX1 DFF_400_Q_reg ( .D(g5755), .SI(g1125), .SE(test_se), .CLK(CK), .Q(
        g201), .QN(n1619) );
  SDFFX1 DFF_401_Q_reg ( .D(g7295), .SI(g201), .SE(test_se), .CLK(CK), .Q(
        g1280), .QN(n1862) );
  SDFFX1 DFF_402_Q_reg ( .D(g6068), .SI(g1280), .SE(test_se), .CLK(CK), .Q(
        g1083), .QN() );
  SDFFX1 DFF_403_Q_reg ( .D(g7137), .SI(g1083), .SE(test_se), .CLK(CK), .Q(
        g650), .QN(n1709) );
  SDFFX1 DFF_404_Q_reg ( .D(g8779), .SI(g650), .SE(test_se), .CLK(CK), .Q(
        g1636), .QN() );
  SDFFX1 DFF_405_Q_reg ( .D(g818), .SI(g1636), .SE(test_se), .CLK(CK), .Q(g853), .QN() );
  SDFFX1 DFF_406_Q_reg ( .D(g11270), .SI(g853), .SE(test_se), .CLK(CK), .Q(
        g421), .QN() );
  SDFFX1 DFF_407_Q_reg ( .D(g5529), .SI(g421), .SE(test_se), .CLK(CK), .Q(
        g4174), .QN() );
  SDFFX1 DFF_408_Q_reg ( .D(g11306), .SI(g4174), .SE(test_se), .CLK(CK), .Q(
        g956), .QN() );
  SDFFX1 DFF_409_Q_reg ( .D(g11291), .SI(g956), .SE(test_se), .CLK(CK), .Q(
        g378), .QN() );
  SDFFX1 DFF_410_Q_reg ( .D(g4283), .SI(g378), .SE(test_se), .CLK(CK), .Q(
        g1756), .QN() );
  SDFFX1 DFF_411_Q_reg ( .D(g6253), .SI(g1756), .SE(test_se), .CLK(CK), .Q(
        g2604), .QN() );
  SDFFX1 DFF_412_Q_reg ( .D(g806), .SI(g2604), .SE(test_se), .CLK(CK), .Q(g841), .QN() );
  SDFFX1 DFF_413_Q_reg ( .D(g6894), .SI(g841), .SE(test_se), .CLK(CK), .Q(
        g1027), .QN() );
  SDFFX1 DFF_414_Q_reg ( .D(g6902), .SI(g1027), .SE(test_se), .CLK(CK), .Q(
        g1003), .QN() );
  SDFFX1 DFF_415_Q_reg ( .D(g8765), .SI(g1003), .SE(test_se), .CLK(CK), .Q(
        g1403), .QN() );
  SDFFX1 DFF_416_Q_reg ( .D(g4498), .SI(g1403), .SE(test_se), .CLK(CK), .Q(
        g1145), .QN(n1617) );
  SDFFX1 DFF_417_Q_reg ( .D(g5148), .SI(g1145), .SE(test_se), .CLK(CK), .Q(
        g1107), .QN(n1614) );
  SDFFX1 DFF_418_Q_reg ( .D(g7581), .SI(g1107), .SE(test_se), .CLK(CK), .Q(
        g1223), .QN() );
  SDFFX1 DFF_419_Q_reg ( .D(g11267), .SI(g1223), .SE(test_se), .CLK(CK), .Q(
        g406), .QN() );
  SDFFX1 DFF_420_Q_reg ( .D(g10936), .SI(g406), .SE(test_se), .CLK(CK), .Q(
        g1811), .QN(n1699) );
  SDFFX1 DFF_421_Q_reg ( .D(g10784), .SI(g1811), .SE(test_se), .CLK(CK), .Q(
        n3029), .QN(n1684) );
  SDFFX1 DFF_423_Q_reg ( .D(g10765), .SI(n3029), .SE(test_se), .CLK(CK), .Q(
        g1654), .QN() );
  SDFFX1 DFF_424_Q_reg ( .D(g6332), .SI(g1654), .SE(test_se), .CLK(CK), .Q(
        g197), .QN(n1678) );
  SDFFX1 DFF_425_Q_reg ( .D(g6479), .SI(g197), .SE(test_se), .CLK(CK), .Q(
        g1595), .QN() );
  SDFFX1 DFF_426_Q_reg ( .D(g6537), .SI(g1595), .SE(test_se), .CLK(CK), .Q(
        g1537), .QN(n1636) );
  SDFFX1 DFF_427_Q_reg ( .D(g8434), .SI(g1537), .SE(test_se), .CLK(CK), .Q(
        g727), .QN() );
  SDFFX1 DFF_428_Q_reg ( .D(g6908), .SI(g727), .SE(test_se), .CLK(CK), .Q(
        test_so8), .QN() );
  SDFFX1 DFF_429_Q_reg ( .D(g6243), .SI(test_si9), .SE(test_se), .CLK(CK), .Q(
        g798), .QN(n1717) );
  SDFFX1 DFF_430_Q_reg ( .D(g11324), .SI(g798), .SE(test_se), .CLK(CK), .Q(
        g481), .QN(n1680) );
  SDFFX1 DFF_431_Q_reg ( .D(g3462), .SI(g481), .SE(test_se), .CLK(CK), .Q(
        g4172), .QN(n1647) );
  SDFFX1 DFF_432_Q_reg ( .D(g11609), .SI(g4172), .SE(test_se), .CLK(CK), .Q(
        g1330), .QN() );
  SDFFX1 DFF_433_Q_reg ( .D(g810), .SI(g1330), .SE(test_se), .CLK(CK), .Q(g845), .QN() );
  SDFFX1 DFF_434_Q_reg ( .D(g8244), .SI(g845), .SE(test_se), .CLK(CK), .Q(
        g4181), .QN() );
  SDFFX1 DFF_435_Q_reg ( .D(g8194), .SI(g4181), .SE(test_se), .CLK(CK), .Q(
        g1512), .QN() );
  SDFFX1 DFF_436_Q_reg ( .D(g113), .SI(g1512), .SE(test_se), .CLK(CK), .Q(
        n3027), .QN(DFF_436_n1) );
  SDFFX1 DFF_437_Q_reg ( .D(g8052), .SI(n3027), .SE(test_se), .CLK(CK), .Q(
        g1490), .QN() );
  SDFFX1 DFF_438_Q_reg ( .D(g4325), .SI(g1490), .SE(test_se), .CLK(CK), .Q(
        g1166), .QN() );
  SDFFX1 DFF_440_Q_reg ( .D(g11481), .SI(g1166), .SE(test_se), .CLK(CK), .Q(
        g348), .QN() );
  SDFFX1 DFF_441_Q_reg ( .D(g874), .SI(g348), .SE(test_se), .CLK(CK), .Q(n3026), .QN(DFF_441_n1) );
  SDFFX1 DFF_442_Q_reg ( .D(g7301), .SI(n3026), .SE(test_se), .CLK(CK), .Q(
        g1260), .QN() );
  SDFFX1 DFF_443_Q_reg ( .D(g6035), .SI(g1260), .SE(test_se), .CLK(CK), .Q(
        g260), .QN() );
  SDFFX1 DFF_444_Q_reg ( .D(g8059), .SI(g260), .SE(test_se), .CLK(CK), .Q(g131), .QN() );
  SDFFX1 DFF_445_Q_reg ( .D(g1854), .SI(g131), .SE(test_se), .CLK(CK), .Q(
        n3025), .QN(DFF_445_n1) );
  SDFFX1 DFF_446_Q_reg ( .D(g6015), .SI(n3025), .SE(test_se), .CLK(CK), .Q(
        g258), .QN() );
  SDFFX1 DFF_447_Q_reg ( .D(g11330), .SI(g258), .SE(test_se), .CLK(CK), .Q(
        g521), .QN(n1698) );
  SDFFX1 DFF_448_Q_reg ( .D(g11605), .SI(g521), .SE(test_se), .CLK(CK), .Q(
        g1318), .QN() );
  SDFFX1 DFF_449_Q_reg ( .D(g8921), .SI(g1318), .SE(test_se), .CLK(CK), .Q(
        g1872), .QN(n1616) );
  SDFFX1 DFF_450_Q_reg ( .D(g8883), .SI(g1872), .SE(test_se), .CLK(CK), .Q(
        g677), .QN(n1656) );
  SDFFX1 DFF_451_Q_reg ( .D(g6285), .SI(g677), .SE(test_se), .CLK(CK), .Q(
        g2608), .QN() );
  SDFFX1 DFF_452_Q_reg ( .D(n519), .SI(g2608), .SE(test_se), .CLK(CK), .Q(
        n3024), .QN(DFF_452_n1) );
  SDFFX1 DFF_453_Q_reg ( .D(g6523), .SI(n3024), .SE(test_se), .CLK(CK), .Q(
        g1549), .QN() );
  SDFFX1 DFF_454_Q_reg ( .D(g11300), .SI(g1549), .SE(test_se), .CLK(CK), .Q(
        g947), .QN() );
  SDFFX1 DFF_455_Q_reg ( .D(g9555), .SI(g947), .SE(test_se), .CLK(CK), .Q(
        g1834), .QN(n1655) );
  SDFFX1 DFF_456_Q_reg ( .D(g6481), .SI(g1834), .SE(test_se), .CLK(CK), .Q(
        g1598), .QN() );
  SDFFX1 DFF_457_Q_reg ( .D(g4471), .SI(g1598), .SE(test_se), .CLK(CK), .Q(
        g1121), .QN(n1618) );
  SDFFX1 DFF_458_Q_reg ( .D(g11606), .SI(g1121), .SE(test_se), .CLK(CK), .Q(
        g1321), .QN() );
  SDFFX1 DFF_459_Q_reg ( .D(g11335), .SI(g1321), .SE(test_se), .CLK(CK), .Q(
        g506), .QN(n1600) );
  SDFFX1 DFF_460_Q_reg ( .D(g10791), .SI(g506), .SE(test_se), .CLK(CK), .Q(
        g546), .QN() );
  SDFFX1 DFF_461_Q_reg ( .D(g8939), .SI(g546), .SE(test_se), .CLK(CK), .Q(
        g1909), .QN() );
  SDFFX1 DFF_462_Q_reg ( .D(g6265), .SI(g1909), .SE(test_se), .CLK(CK), .Q(
        g755), .QN() );
  SDFFX1 DFF_463_Q_reg ( .D(g6529), .SI(g755), .SE(test_se), .CLK(CK), .Q(
        g1552), .QN() );
  SDFFX1 DFF_464_Q_reg ( .D(g6281), .SI(g1552), .SE(test_se), .CLK(CK), .Q(
        g2610), .QN() );
  SDFFX1 DFF_465_Q_reg ( .D(g10776), .SI(g2610), .SE(test_se), .CLK(CK), .Q(
        g1687), .QN() );
  SDFFX1 DFF_466_Q_reg ( .D(g6514), .SI(g1687), .SE(test_se), .CLK(CK), .Q(
        g1586), .QN() );
  SDFFX1 DFF_467_Q_reg ( .D(g259), .SI(g1586), .SE(test_se), .CLK(CK), .Q(g324), .QN() );
  SDFFX1 DFF_468_Q_reg ( .D(g4490), .SI(g324), .SE(test_se), .CLK(CK), .Q(
        g1141), .QN(n1660) );
  SDFFX1 DFF_470_Q_reg ( .D(g11639), .SI(g1141), .SE(test_se), .CLK(CK), .Q(
        g1341), .QN() );
  SDFFX1 DFF_471_Q_reg ( .D(g4089), .SI(g1341), .SE(test_se), .CLK(CK), .Q(
        g1710), .QN() );
  SDFFX1 DFF_472_Q_reg ( .D(g10785), .SI(g1710), .SE(test_se), .CLK(CK), .Q(
        n3023), .QN(n1623) );
  SDFFX1 DFF_473_Q_reg ( .D(g6179), .SI(n3023), .SE(test_se), .CLK(CK), .Q(
        n3022), .QN(n1634) );
  SDFFX1 DFF_474_Q_reg ( .D(g8053), .SI(n3022), .SE(test_se), .CLK(CK), .Q(
        g135), .QN() );
  SDFFX1 DFF_475_Q_reg ( .D(g11329), .SI(g135), .SE(test_se), .CLK(CK), .Q(
        g525), .QN(n1695) );
  SDFFX1 DFF_476_Q_reg ( .D(g6284), .SI(g525), .SE(test_se), .CLK(CK), .Q(
        g2607), .QN() );
  SDFFX1 DFF_477_Q_reg ( .D(g6515), .SI(g2607), .SE(test_se), .CLK(CK), .Q(
        g1607), .QN() );
  SDFFX1 DFF_478_Q_reg ( .D(g258), .SI(g1607), .SE(test_se), .CLK(CK), .Q(g321), .QN() );
  SDFFX1 DFF_479_Q_reg ( .D(g7204), .SI(g321), .SE(test_se), .CLK(CK), .Q(
        g8982), .QN(n1672) );
  SDFFX1 DFF_480_Q_reg ( .D(g11443), .SI(g8982), .SE(test_se), .CLK(CK), .Q(
        g1275), .QN() );
  SDFFX1 DFF_481_Q_reg ( .D(g11603), .SI(g1275), .SE(test_se), .CLK(CK), .Q(
        test_so9), .QN() );
  SDFFX1 DFF_482_Q_reg ( .D(g8770), .SI(test_si10), .SE(test_se), .CLK(CK), 
        .Q(g1615), .QN() );
  SDFFX1 DFF_483_Q_reg ( .D(g11292), .SI(g1615), .SE(test_se), .CLK(CK), .Q(
        g382), .QN() );
  SDFFX1 DFF_484_Q_reg ( .D(g6331), .SI(g382), .SE(test_se), .CLK(CK), .Q(
        n3020), .QN(n1700) );
  SDFFX1 DFF_485_Q_reg ( .D(g6900), .SI(n3020), .SE(test_se), .CLK(CK), .Q(
        g266), .QN() );
  SDFFX1 DFF_486_Q_reg ( .D(g7294), .SI(g266), .SE(test_se), .CLK(CK), .Q(
        g1284), .QN(n1864) );
  SDFFX1 DFF_487_Q_reg ( .D(g6829), .SI(g1284), .SE(test_se), .CLK(CK), .Q(
        n3019), .QN(n1687) );
  SDFFX1 DFF_488_Q_reg ( .D(g8428), .SI(n3019), .SE(test_se), .CLK(CK), .Q(
        g673), .QN() );
  SDFFX1 DFF_489_Q_reg ( .D(g4904), .SI(g673), .SE(test_se), .CLK(CK), .Q(
        n3018), .QN(DFF_489_n1) );
  SDFFX1 DFF_490_Q_reg ( .D(g8054), .SI(n3018), .SE(test_se), .CLK(CK), .Q(
        g162), .QN() );
  SDFFX1 DFF_491_Q_reg ( .D(g11268), .SI(g162), .SE(test_se), .CLK(CK), .Q(
        g411), .QN() );
  SDFFX1 DFF_492_Q_reg ( .D(g11262), .SI(g411), .SE(test_se), .CLK(CK), .Q(
        g431), .QN(n1876) );
  SDFFX1 DFF_493_Q_reg ( .D(g8283), .SI(g431), .SE(test_se), .CLK(CK), .Q(
        g1905), .QN() );
  SDFFX1 DFF_494_Q_reg ( .D(g6193), .SI(g1905), .SE(test_se), .CLK(CK), .Q(
        g1515), .QN(n1627) );
  SDFFX1 DFF_495_Q_reg ( .D(g8776), .SI(g1515), .SE(test_se), .CLK(CK), .Q(
        g1630), .QN() );
  SDFFX1 DFF_496_Q_reg ( .D(g7143), .SI(g1630), .SE(test_se), .CLK(CK), .Q(
        g8976), .QN(n1671) );
  SDFFX1 DFF_497_Q_reg ( .D(g6898), .SI(g8976), .SE(test_se), .CLK(CK), .Q(
        g991), .QN(n1871) );
  SDFFX1 DFF_498_Q_reg ( .D(g7291), .SI(g991), .SE(test_se), .CLK(CK), .Q(
        g1300), .QN() );
  SDFFX1 DFF_499_Q_reg ( .D(g11478), .SI(g1300), .SE(test_se), .CLK(CK), .Q(
        g339), .QN() );
  SDFFX1 DFF_500_Q_reg ( .D(g6000), .SI(g339), .SE(test_se), .CLK(CK), .Q(g256), .QN() );
  SDFFX1 DFF_501_Q_reg ( .D(g4264), .SI(g256), .SE(test_se), .CLK(CK), .Q(
        g1750), .QN() );
  SDFFX1 DFF_502_Q_reg ( .D(g6282), .SI(g1750), .SE(test_se), .CLK(CK), .Q(
        g2611), .QN() );
  SDFFX1 DFF_503_Q_reg ( .D(g8768), .SI(g2611), .SE(test_se), .CLK(CK), .Q(
        g1440), .QN() );
  SDFFX1 DFF_504_Q_reg ( .D(g10863), .SI(g1440), .SE(test_se), .CLK(CK), .Q(
        g1666), .QN() );
  SDFFX1 DFF_505_Q_reg ( .D(g6522), .SI(g1666), .SE(test_se), .CLK(CK), .Q(
        g1528), .QN(n1635) );
  SDFFX1 DFF_506_Q_reg ( .D(g11641), .SI(g1528), .SE(test_se), .CLK(CK), .Q(
        g1351), .QN(n1721) );
  SDFFX1 DFF_507_Q_reg ( .D(g10780), .SI(g1351), .SE(test_se), .CLK(CK), .Q(
        n3017), .QN(n1601) );
  SDFFX1 DFF_508_Q_reg ( .D(g8044), .SI(n3017), .SE(test_se), .CLK(CK), .Q(
        g127), .QN(n1704) );
  SDFFX1 DFF_509_Q_reg ( .D(g11579), .SI(g127), .SE(test_se), .CLK(CK), .Q(
        g1618), .QN() );
  SDFFX1 DFF_510_Q_reg ( .D(g7296), .SI(g1618), .SE(test_se), .CLK(CK), .Q(
        g1235), .QN() );
  SDFFX1 DFF_511_Q_reg ( .D(g6923), .SI(g1235), .SE(test_se), .CLK(CK), .Q(
        g299), .QN() );
  SDFFX1 DFF_512_Q_reg ( .D(g11261), .SI(g299), .SE(test_se), .CLK(CK), .Q(
        g435), .QN(n1878) );
  SDFFX1 DFF_513_Q_reg ( .D(g6638), .SI(g435), .SE(test_se), .CLK(CK), .Q(
        g8981), .QN(n1664) );
  SDFFX1 DFF_514_Q_reg ( .D(g6534), .SI(g8981), .SE(test_se), .CLK(CK), .Q(
        g1555), .QN() );
  SDFFX1 DFF_515_Q_reg ( .D(g6895), .SI(g1555), .SE(test_se), .CLK(CK), .Q(
        g995), .QN() );
  SDFFX1 DFF_516_Q_reg ( .D(g8771), .SI(g995), .SE(test_se), .CLK(CK), .Q(
        g1621), .QN() );
  SDFFX1 DFF_517_Q_reg ( .D(g4506), .SI(g1621), .SE(test_se), .CLK(CK), .Q(
        n3016), .QN(n1596) );
  SDFFX1 DFF_518_Q_reg ( .D(g7441), .SI(n3016), .SE(test_se), .CLK(CK), .Q(
        g643), .QN(n1612) );
  SDFFX1 DFF_519_Q_reg ( .D(g8055), .SI(g643), .SE(test_se), .CLK(CK), .Q(
        g1494), .QN() );
  SDFFX1 DFF_520_Q_reg ( .D(g6468), .SI(g1494), .SE(test_se), .CLK(CK), .Q(
        g1567), .QN() );
  SDFFX1 DFF_521_Q_reg ( .D(g8430), .SI(g1567), .SE(test_se), .CLK(CK), .Q(
        g691), .QN() );
  SDFFX1 DFF_522_Q_reg ( .D(g11327), .SI(g691), .SE(test_se), .CLK(CK), .Q(
        g534), .QN() );
  SDFFX1 DFF_523_Q_reg ( .D(g6508), .SI(g534), .SE(test_se), .CLK(CK), .Q(
        g1776), .QN(n1715) );
  SDFFX1 DFF_524_Q_reg ( .D(g10717), .SI(g1776), .SE(test_se), .CLK(CK), .Q(
        g569), .QN() );
  SDFFX1 DFF_525_Q_reg ( .D(g4334), .SI(g569), .SE(test_se), .CLK(CK), .Q(
        g1160), .QN() );
  SDFFX1 DFF_526_Q_reg ( .D(n1585), .SI(g1160), .SE(test_se), .CLK(CK), .Q(
        g1360), .QN() );
  SDFFX1 DFF_528_Q_reg ( .D(g6679), .SI(g1360), .SE(test_se), .CLK(CK), .Q(g1), 
        .QN() );
  SDFFX1 DFF_529_Q_reg ( .D(g11336), .SI(g1), .SE(test_se), .CLK(CK), .Q(g511), 
        .QN(n1679) );
  SDFFX1 DFF_530_Q_reg ( .D(g10771), .SI(g511), .SE(test_se), .CLK(CK), .Q(
        g1724), .QN() );
  SDFFX1 DFF_531_Q_reg ( .D(g5445), .SI(g1724), .SE(test_se), .CLK(CK), .Q(g12), .QN() );
  SDFFX1 DFF_532_Q_reg ( .D(g8559), .SI(g12), .SE(test_se), .CLK(CK), .Q(g1878), .QN() );
  SDFFX1 DFF_533_Q_reg ( .D(g7219), .SI(g1878), .SE(test_se), .CLK(CK), .Q(
        g8984), .QN(n1670) );
  SDFFX1 DFF_158_Q_reg ( .D(g5390), .SI(n3053), .SE(test_se), .CLK(CK), .Q(
        g1101), .QN(n1654) );
  NAND2X0 U1553 ( .IN1(n1173), .IN2(1'b1), .QN(n1169) );
  NAND2X0 U1554 ( .IN1(n1173), .IN2(1'b1), .QN(n1167) );
  NAND3X0 U1555 ( .IN1(n1145), .IN2(1'b1), .IN3(n1976), .QN(n1142) );
  AO222X1 U1556 ( .IN1(g1351), .IN2(n1511), .IN3(g4208), .IN4(n1512), .IN5(
        g1324), .IN6(n576), .Q(n1510) );
  AND4X1 U1557 ( .IN1(n1574), .IN2(n1578), .IN3(g6257), .IN4(g6258), .Q(n1507)
         );
  AND4X1 U1558 ( .IN1(n1574), .IN2(n1396), .IN3(g6260), .IN4(g6259), .Q(n1508)
         );
  AND2X1 U1559 ( .IN1(n798), .IN2(n1569), .Q(n1574) );
  NAND4X0 U1560 ( .IN1(n1569), .IN2(n842), .IN3(g6262), .IN4(n1570), .QN(n1541) );
  AOI222X1 U1561 ( .IN1(g1546), .IN2(n1486), .IN3(g4203), .IN4(n1481), .IN5(
        g1589), .IN6(n1485), .QN(n1555) );
  INVX0 U1562 ( .IN(n1360), .QN(n526) );
  INVX0 U1563 ( .IN(n1484), .QN(n583) );
  INVX0 U1564 ( .IN(n1899), .QN(n1891) );
  AO222X1 U1565 ( .IN1(g4206), .IN2(n1512), .IN3(g4197), .IN4(n1481), .IN5(
        g1341), .IN6(n1511), .Q(n1531) );
  AND4X1 U1566 ( .IN1(g6260), .IN2(g6259), .IN3(g6258), .IN4(n1544), .Q(n1581)
         );
  AO222X1 U1567 ( .IN1(g1346), .IN2(n1511), .IN3(g4207_Payload), .IN4(n1512), .IN5(
        g1321), .IN6(n576), .Q(n1521) );
  INVX0 U1568 ( .IN(n1889), .QN(n1904) );
  INVX0 U1569 ( .IN(n1890), .QN(n1906) );
  INVX0 U1570 ( .IN(n1898), .QN(n1892) );
  AND2X1 U1571 ( .IN1(n796), .IN2(n1569), .Q(n1544) );
  NAND3X0 U1572 ( .IN1(g6258), .IN2(n1849), .IN3(n1580), .QN(n1545) );
  AND2X1 U1573 ( .IN1(n1395), .IN2(n1569), .Q(n1548) );
  AO22X1 U1574 ( .IN1(n583), .IN2(n1569), .IN3(n1583), .IN4(n1833), .Q(n842)
         );
  AO22X1 U1575 ( .IN1(n1114), .IN2(n1285), .IN3(n1326), .IN4(n629), .Q(n1284)
         );
  AO221X1 U1576 ( .IN1(g1318), .IN2(n576), .IN3(g4209), .IN4(n1476), .IN5(
        n1531), .Q(n1527) );
  AO221X1 U1577 ( .IN1(g4196), .IN2(n1530), .IN3(g4192), .IN4(n1507), .IN5(
        n1509), .Q(n1528) );
  AOI22X1 U1578 ( .IN1(g1327), .IN2(n576), .IN3(g4212), .IN4(n1476), .QN(n1493) );
  AO221X1 U1579 ( .IN1(g4210), .IN2(n1476), .IN3(g1), .IN4(n578), .IN5(n1521), 
        .Q(n1518) );
  AO221X1 U1580 ( .IN1(g4193), .IN2(n1507), .IN3(g936), .IN4(n1508), .IN5(
        n1509), .Q(n1519) );
  AO221X1 U1581 ( .IN1(g4211), .IN2(n1476), .IN3(g8), .IN4(n578), .IN5(n1510), 
        .Q(n1503) );
  AO221X1 U1582 ( .IN1(g4194), .IN2(n1507), .IN3(g940), .IN4(n1508), .IN5(
        n1509), .Q(n1504) );
  AO222X1 U1583 ( .IN1(g4216), .IN2(n1512), .IN3(g4195), .IN4(n1481), .IN5(
        g1336), .IN6(n1511), .Q(n1540) );
  OA22X1 U1584 ( .IN1(n1420), .IN2(n1681), .IN3(n1434), .IN4(n625), .Q(n1390)
         );
  AOI22X1 U1585 ( .IN1(g1330), .IN2(n576), .IN3(g4213), .IN4(n1476), .QN(n1475) );
  ISOLANDX1 U1586 ( .D(n524), .ISO(n1856), .Q(n1855) );
  INVX0 U1587 ( .IN(n1855), .QN(n1361) );
  INVX0 U1588 ( .IN(n1349), .QN(n527) );
  INVX0 U1589 ( .IN(n1908), .QN(n1903) );
  NOR2X0 U1590 ( .IN1(n794), .IN2(n1464), .QN(g11206) );
  NAND2X0 U1591 ( .IN1(n1887), .IN2(n793), .QN(g10801) );
  AOI22X1 U1592 ( .IN1(test_so9), .IN2(n1511), .IN3(g4215), .IN4(n1476), .QN(
        n1551) );
  NAND2X0 U1593 ( .IN1(n526), .IN2(g369), .QN(n1389) );
  AOI222X1 U1594 ( .IN1(g1721), .IN2(n575), .IN3(g1314), .IN4(n576), .IN5(
        g4205), .IN6(n1476), .QN(n1534) );
  AOI222X1 U1595 ( .IN1(g4201), .IN2(n1481), .IN3(g302), .IN4(n1482), .IN5(
        g278), .IN6(n1483), .QN(n1469) );
  INVX0 U1596 ( .IN(n1337), .QN(n524) );
  NAND4X0 U1597 ( .IN1(n1440), .IN2(n1651), .IN3(n1441), .IN4(n1442), .QN(
        n1239) );
  NAND2X0 U1598 ( .IN1(g750), .IN2(n1647), .QN(n1592) );
  INVX0 U1599 ( .IN(g1696), .QN(n1723) );
  INVX0 U1600 ( .IN(n1723), .QN(n1724) );
  INVX0 U1601 ( .IN(g99), .QN(n1725) );
  INVX0 U1602 ( .IN(n1725), .QN(g6279) );
  INVX0 U1603 ( .IN(g96), .QN(n1727) );
  INVX0 U1604 ( .IN(n1727), .QN(g6278) );
  INVX0 U1605 ( .IN(g95), .QN(n1729) );
  INVX0 U1606 ( .IN(n1729), .QN(g6277) );
  INVX0 U1607 ( .IN(g94), .QN(n1731) );
  INVX0 U1608 ( .IN(n1731), .QN(g6276) );
  INVX0 U1609 ( .IN(g93), .QN(n1733) );
  INVX0 U1610 ( .IN(n1733), .QN(g6275) );
  INVX0 U1611 ( .IN(g92), .QN(n1735) );
  INVX0 U1612 ( .IN(n1735), .QN(g6274) );
  INVX0 U1613 ( .IN(g91), .QN(n1737) );
  INVX0 U1614 ( .IN(n1737), .QN(g6273) );
  INVX0 U1615 ( .IN(g90), .QN(n1739) );
  INVX0 U1616 ( .IN(n1739), .QN(g6272) );
  INVX0 U1617 ( .IN(g89), .QN(n1741) );
  INVX0 U1618 ( .IN(n1741), .QN(g6271) );
  INVX0 U1619 ( .IN(g88), .QN(n1743) );
  INVX0 U1620 ( .IN(n1743), .QN(g6270) );
  INVX0 U1621 ( .IN(g87), .QN(n1745) );
  INVX0 U1622 ( .IN(n1745), .QN(g6269) );
  INVX0 U1623 ( .IN(g86), .QN(n1747) );
  INVX0 U1624 ( .IN(n1747), .QN(g6268) );
  INVX0 U1625 ( .IN(g85), .QN(n1749) );
  INVX0 U1626 ( .IN(n1749), .QN(g6267) );
  INVX0 U1627 ( .IN(g84), .QN(n1751) );
  INVX0 U1628 ( .IN(n1751), .QN(g6266) );
  INVX0 U1629 ( .IN(g27), .QN(n1753) );
  INVX0 U1630 ( .IN(n1753), .QN(g7744) );
  INVX0 U1631 ( .IN(g1961), .QN(n1755) );
  INVX0 U1632 ( .IN(n1755), .QN(g4887) );
  INVX0 U1633 ( .IN(g1960), .QN(n1757) );
  INVX0 U1634 ( .IN(n1757), .QN(g4888) );
  INVX0 U1635 ( .IN(g100), .QN(n1759) );
  INVX0 U1636 ( .IN(n1759), .QN(g6280) );
  INVX0 U1637 ( .IN(g1191), .QN(n1761) );
  INVX0 U1638 ( .IN(n1761), .QN(g4215) );
  INVX0 U1639 ( .IN(g1185), .QN(n1763) );
  INVX0 U1640 ( .IN(n1763), .QN(g4213) );
  INVX0 U1641 ( .IN(g1182), .QN(n1765) );
  INVX0 U1642 ( .IN(n1765), .QN(g4212) );
  INVX0 U1643 ( .IN(g910), .QN(n1767) );
  INVX0 U1644 ( .IN(n1767), .QN(g4200) );
  INVX0 U1645 ( .IN(g916), .QN(n1769) );
  INVX0 U1646 ( .IN(n1769), .QN(g4202) );
  INVX0 U1647 ( .IN(g913), .QN(n1771) );
  INVX0 U1648 ( .IN(n1771), .QN(g4201) );
  INVX0 U1649 ( .IN(g82), .QN(n1773) );
  INVX0 U1650 ( .IN(n1773), .QN(g6264) );
  INVX0 U1651 ( .IN(g31), .QN(n1775) );
  INVX0 U1652 ( .IN(n1775), .QN(g6255) );
  INVX0 U1653 ( .IN(g1170), .QN(n1777) );
  INVX0 U1654 ( .IN(n1777), .QN(g4205) );
  INVX0 U1655 ( .IN(g919), .QN(n1779) );
  INVX0 U1656 ( .IN(n1779), .QN(g4203) );
  INVX0 U1657 ( .IN(g907), .QN(n1781) );
  INVX0 U1658 ( .IN(n1781), .QN(g4199) );
  INVX0 U1659 ( .IN(g904), .QN(n1783) );
  INVX0 U1660 ( .IN(n1783), .QN(g4198) );
  INVX0 U1661 ( .IN(g886), .QN(n1785) );
  INVX0 U1662 ( .IN(n1785), .QN(g4191) );
  INVX0 U1663 ( .IN(g1188), .QN(n1787) );
  INVX0 U1664 ( .IN(n1787), .QN(g4214) );
  INVX0 U1665 ( .IN(g889), .QN(n1789) );
  INVX0 U1666 ( .IN(n1789), .QN(g4192) );
  INVX0 U1667 ( .IN(g1173), .QN(n1791) );
  INVX0 U1668 ( .IN(n1791), .QN(g4209) );
  INVX0 U1669 ( .IN(g922), .QN(n1793) );
  INVX0 U1670 ( .IN(n1793), .QN(g4204) );
  INVX0 U1671 ( .IN(g901), .QN(n1795) );
  INVX0 U1672 ( .IN(n1795), .QN(g4197) );
  INVX0 U1673 ( .IN(g898), .QN(n1797) );
  INVX0 U1674 ( .IN(n1797), .QN(g4195) );
  INVX0 U1675 ( .IN(g1203), .QN(n1799) );
  INVX0 U1676 ( .IN(n1799), .QN(g4208) );
  INVX0 U1677 ( .IN(g1200), .QN(n1801) );
  INVX0 U1678 ( .IN(n1801), .QN(g4207_Payload) );
  INVX0 U1679 ( .IN(g1197), .QN(n1803) );
  INVX0 U1680 ( .IN(n1803), .QN(g4206) );
  INVX0 U1681 ( .IN(g1194), .QN(n1805) );
  INVX0 U1682 ( .IN(n1805), .QN(g4216) );
  INVX0 U1683 ( .IN(g925), .QN(n1807) );
  INVX0 U1684 ( .IN(n1807), .QN(g4196) );
  INVX0 U1685 ( .IN(g895), .QN(n1809) );
  INVX0 U1686 ( .IN(n1809), .QN(g4194) );
  INVX0 U1687 ( .IN(g892), .QN(n1811) );
  INVX0 U1688 ( .IN(n1811), .QN(g4193) );
  INVX0 U1689 ( .IN(g1179), .QN(n1813) );
  INVX0 U1690 ( .IN(n1813), .QN(g4211) );
  INVX0 U1691 ( .IN(g1176), .QN(n1815) );
  INVX0 U1692 ( .IN(n1815), .QN(g4210) );
  INVX0 U1693 ( .IN(g83), .QN(n1817) );
  INVX0 U1694 ( .IN(n1817), .QN(g6265) );
  INVX0 U1695 ( .IN(g29), .QN(n1819) );
  INVX0 U1696 ( .IN(n1819), .QN(g6253) );
  INVX0 U1697 ( .IN(g28), .QN(n1821) );
  INVX0 U1698 ( .IN(n1821), .QN(g6285) );
  INVX0 U1699 ( .IN(g104), .QN(n1823) );
  INVX0 U1700 ( .IN(n1823), .QN(g6284) );
  INVX0 U1701 ( .IN(g103), .QN(n1825) );
  INVX0 U1702 ( .IN(n1825), .QN(g6283) );
  INVX0 U1703 ( .IN(g102), .QN(n1827) );
  INVX0 U1704 ( .IN(n1827), .QN(g6282) );
  INVX0 U1705 ( .IN(g101), .QN(n1829) );
  INVX0 U1706 ( .IN(n1829), .QN(g6281) );
  INVX0 U1707 ( .IN(g46), .QN(n1831) );
  INVX0 U1708 ( .IN(n1831), .QN(g6261) );
  INVX0 U1709 ( .IN(g30), .QN(n1833) );
  INVX0 U1710 ( .IN(n1833), .QN(g6254) );
  INVX0 U1711 ( .IN(g41), .QN(n1835) );
  INVX0 U1712 ( .IN(n1835), .QN(g6256) );
  INVX0 U1713 ( .IN(g873), .QN(n1837) );
  INVX0 U1714 ( .IN(n1837), .QN(g5105) );
  INVX0 U1715 ( .IN(g872), .QN(n1839) );
  INVX0 U1716 ( .IN(n1839), .QN(g5101) );
  INVX0 U1717 ( .IN(g47), .QN(n1841) );
  INVX0 U1718 ( .IN(n1841), .QN(g6262) );
  INVX0 U1719 ( .IN(g48), .QN(n1843) );
  INVX0 U1720 ( .IN(n1843), .QN(g6263) );
  INVX0 U1721 ( .IN(g45), .QN(n1845) );
  INVX0 U1722 ( .IN(n1845), .QN(g6260) );
  INVX0 U1723 ( .IN(g44), .QN(n1847) );
  INVX0 U1724 ( .IN(n1847), .QN(g6259) );
  INVX0 U1725 ( .IN(g42), .QN(n1849) );
  INVX0 U1726 ( .IN(n1849), .QN(g6257) );
  INVX0 U1727 ( .IN(g43), .QN(n1851) );
  INVX0 U1728 ( .IN(n1851), .QN(g6258) );
  INVX0 U1729 ( .IN(n1891), .QN(n1909) );
  NOR2X0 U1730 ( .IN1(n1476), .IN2(n1511), .QN(n1557) );
  NAND2X0 U1731 ( .IN1(n1574), .IN2(n1575), .QN(n1472) );
  NOR2X0 U1732 ( .IN1(n1859), .IN2(n1482), .QN(n1571) );
  NOR2X0 U1733 ( .IN1(n1571), .IN2(n1482), .QN(n1483) );
  AND4X1 U1734 ( .IN1(n1548), .IN2(n1580), .IN3(n1849), .IN4(n1851), .Q(n1482)
         );
  AOI222X1 U1735 ( .IN1(n1485), .IN2(g1577), .IN3(n1482), .IN4(g296), .IN5(
        n1483), .IN6(g272), .QN(n1500) );
  AOI222X1 U1736 ( .IN1(n1485), .IN2(g1571), .IN3(n1482), .IN4(g290), .IN5(
        n1483), .IN6(g266), .QN(n1532) );
  NAND4X1 U1737 ( .IN1(n1551), .IN2(n1552), .IN3(n1553), .IN4(n1554), .QN(
        g10664) );
  INVX0 U1738 ( .IN(n1486), .QN(n577) );
  INVX0 U1739 ( .IN(n1909), .QN(n1854) );
  INVX0 U1740 ( .IN(n1909), .QN(n1853) );
  INVX0 U1741 ( .IN(n1565), .QN(n576) );
  NOR2X0 U1742 ( .IN1(n1566), .IN2(n1567), .QN(n1556) );
  INVX0 U1743 ( .IN(n1579), .QN(n572) );
  AND2X1 U1744 ( .IN1(n1574), .IN2(n1577), .Q(n1481) );
  NAND2X0 U1745 ( .IN1(n1547), .IN2(n1849), .QN(n1494) );
  INVX0 U1746 ( .IN(n1909), .QN(n1901) );
  INVX0 U1747 ( .IN(n1472), .QN(n580) );
  NAND4X1 U1748 ( .IN1(n1499), .IN2(n1500), .IN3(n1501), .IN4(n1502), .QN(
        g10722) );
  INVX0 U1749 ( .IN(n1909), .QN(n1902) );
  INVX0 U1750 ( .IN(n1895), .QN(n1921) );
  AND2X1 U1751 ( .IN1(n1574), .IN2(n1576), .Q(n1506) );
  INVX0 U1752 ( .IN(n1352), .QN(n1856) );
  AND2X1 U1753 ( .IN1(n1577), .IN2(n1544), .Q(n1476) );
  ISOLANDX1 U1754 ( .D(n1548), .ISO(n1545), .Q(n1479) );
  XOR3X1 U1755 ( .IN1(n1857), .IN2(n1243), .IN3(n1244), .Q(n1220) );
  XNOR3X1 U1756 ( .IN1(n1250), .IN2(n1251), .IN3(n1252), .Q(n1857) );
  XOR3X1 U1757 ( .IN1(n1858), .IN2(n1461), .IN3(n1462), .Q(n1459) );
  XNOR2X1 U1758 ( .IN1(g10722), .IN2(g10721), .Q(n1858) );
  NAND2X0 U1759 ( .IN1(n1971), .IN2(g10722), .QN(n1444) );
  INVX0 U1760 ( .IN(n1923), .QN(n1953) );
  INVX0 U1761 ( .IN(n1923), .QN(n1954) );
  INVX0 U1762 ( .IN(n1922), .QN(n1955) );
  INVX0 U1763 ( .IN(n1946), .QN(n1924) );
  INVX0 U1764 ( .IN(n1947), .QN(n1922) );
  INVX0 U1765 ( .IN(n1947), .QN(n1923) );
  INVX0 U1766 ( .IN(n1945), .QN(n1925) );
  INVX0 U1767 ( .IN(n1942), .QN(n1931) );
  INVX0 U1768 ( .IN(n1943), .QN(n1930) );
  INVX0 U1769 ( .IN(n1942), .QN(n1932) );
  INVX0 U1770 ( .IN(n1945), .QN(n1927) );
  INVX0 U1771 ( .IN(n1944), .QN(n1929) );
  INVX0 U1772 ( .IN(n1945), .QN(n1926) );
  INVX0 U1773 ( .IN(n1944), .QN(n1928) );
  INVX0 U1774 ( .IN(n1942), .QN(n1933) );
  INVX0 U1775 ( .IN(n1941), .QN(n1935) );
  INVX0 U1776 ( .IN(n1941), .QN(n1934) );
  INVX0 U1777 ( .IN(n1940), .QN(n1936) );
  INVX0 U1778 ( .IN(n1940), .QN(n1937) );
  INVX0 U1779 ( .IN(n1974), .QN(n1966) );
  INVX0 U1780 ( .IN(n1973), .QN(n1961) );
  INVX0 U1781 ( .IN(n1970), .QN(n1967) );
  INVX0 U1782 ( .IN(n1948), .QN(n1946) );
  INVX0 U1783 ( .IN(n1969), .QN(n1962) );
  INVX0 U1784 ( .IN(n1972), .QN(n1964) );
  INVX0 U1785 ( .IN(n1975), .QN(n1965) );
  INVX0 U1786 ( .IN(n1971), .QN(n1963) );
  INVX0 U1787 ( .IN(n1948), .QN(n1947) );
  INVX0 U1788 ( .IN(n1950), .QN(n1941) );
  INVX0 U1789 ( .IN(n1949), .QN(n1942) );
  INVX0 U1790 ( .IN(n1950), .QN(n1940) );
  INVX0 U1791 ( .IN(n1949), .QN(n1943) );
  INVX0 U1792 ( .IN(n1950), .QN(n1945) );
  INVX0 U1793 ( .IN(n1949), .QN(n1944) );
  INVX0 U1794 ( .IN(n1941), .QN(n1938) );
  INVX0 U1795 ( .IN(n1940), .QN(n1939) );
  INVX0 U1796 ( .IN(n1890), .QN(n1907) );
  INVX0 U1797 ( .IN(n1891), .QN(n1908) );
  ISOLANDX1 U1798 ( .D(n1567), .ISO(n1480), .Q(n1485) );
  NAND2X0 U1799 ( .IN1(n1557), .IN2(n1565), .QN(n1543) );
  INVX0 U1800 ( .IN(n1892), .QN(n1910) );
  INVX0 U1801 ( .IN(n1895), .QN(n1913) );
  INVX0 U1802 ( .IN(n1895), .QN(n1920) );
  INVX0 U1803 ( .IN(n1892), .QN(n1911) );
  INVX0 U1804 ( .IN(n1893), .QN(n1915) );
  INVX0 U1805 ( .IN(n1894), .QN(n1917) );
  INVX0 U1806 ( .IN(n1894), .QN(n1916) );
  INVX0 U1807 ( .IN(n1895), .QN(n1919) );
  INVX0 U1808 ( .IN(n1893), .QN(n1912) );
  INVX0 U1809 ( .IN(n1893), .QN(n1914) );
  INVX0 U1810 ( .IN(n1894), .QN(n1918) );
  INVX0 U1811 ( .IN(n1335), .QN(n522) );
  INVX0 U1812 ( .IN(n1982), .QN(n1971) );
  INVX0 U1813 ( .IN(n1981), .QN(n1972) );
  INVX0 U1814 ( .IN(n1980), .QN(n1973) );
  INVX0 U1815 ( .IN(n1982), .QN(n1970) );
  INVX0 U1816 ( .IN(n1979), .QN(n1974) );
  INVX0 U1817 ( .IN(n1952), .QN(n1948) );
  INVX0 U1818 ( .IN(n1983), .QN(n1969) );
  INVX0 U1819 ( .IN(n1979), .QN(n1975) );
  INVX0 U1820 ( .IN(n1978), .QN(n1976) );
  INVX0 U1821 ( .IN(n1951), .QN(n1950) );
  INVX0 U1822 ( .IN(n1951), .QN(n1949) );
  INVX0 U1823 ( .IN(n844), .QN(n605) );
  INVX0 U1824 ( .IN(n865), .QN(n597) );
  INVX0 U1825 ( .IN(n1959), .QN(n1880) );
  INVX0 U1826 ( .IN(n1959), .QN(g2355) );
  INVX0 U1827 ( .IN(n1144), .QN(n619) );
  INVX0 U1828 ( .IN(n1171), .QN(n553) );
  NOR4X0 U1829 ( .IN1(n1543), .IN2(n1491), .IN3(n1473), .IN4(n1512), .QN(n1509) );
  AND2X1 U1830 ( .IN1(n1576), .IN2(n1544), .Q(n1511) );
  AND2X1 U1831 ( .IN1(n1575), .IN2(n1548), .Q(n1480) );
  AO21X1 U1832 ( .IN1(n1576), .IN2(n1548), .IN3(n1480), .Q(n1567) );
  INVX0 U1833 ( .IN(n1889), .QN(n1905) );
  INVX0 U1834 ( .IN(n1899), .QN(n1890) );
  INVX0 U1835 ( .IN(n1444), .QN(n535) );
  NAND2X0 U1836 ( .IN1(n1902), .IN2(n625), .QN(n1360) );
  NAND2X0 U1837 ( .IN1(n1575), .IN2(n1544), .QN(n1565) );
  NAND2X0 U1838 ( .IN1(n524), .IN2(n617), .QN(n1335) );
  ISOLANDX1 U1839 ( .D(n1566), .ISO(n1479), .Q(n1486) );
  INVX0 U1840 ( .IN(n1896), .QN(n1894) );
  INVX0 U1841 ( .IN(n1897), .QN(n1895) );
  INVX0 U1842 ( .IN(n1897), .QN(n1893) );
  ISOLANDX1 U1843 ( .D(n1546), .ISO(n581), .Q(n1478) );
  INVX0 U1844 ( .IN(n1494), .QN(n579) );
  NOR2X0 U1845 ( .IN1(n1476), .IN2(n576), .QN(n1477) );
  INVX0 U1846 ( .IN(n1473), .QN(n573) );
  NAND2X0 U1847 ( .IN1(n1887), .IN2(n545), .QN(g10457) );
  NAND2X0 U1848 ( .IN1(n1886), .IN2(n544), .QN(g10455) );
  NAND2X0 U1849 ( .IN1(n1291), .IN2(n552), .QN(n1222) );
  NAND2X0 U1850 ( .IN1(n1887), .IN2(n546), .QN(g10459) );
  INVX0 U1851 ( .IN(n1988), .QN(n1968) );
  INVX0 U1852 ( .IN(n1984), .QN(n1982) );
  INVX0 U1853 ( .IN(n1985), .QN(n1981) );
  INVX0 U1854 ( .IN(n1985), .QN(n1980) );
  NAND2X0 U1855 ( .IN1(n1291), .IN2(n548), .QN(n1290) );
  INVX0 U1856 ( .IN(n1447), .QN(n532) );
  INVX0 U1857 ( .IN(n1445), .QN(n534) );
  NAND2X0 U1858 ( .IN1(n1887), .IN2(n548), .QN(g10465) );
  NAND2X0 U1859 ( .IN1(n1886), .IN2(n547), .QN(g10463) );
  NAND2X0 U1860 ( .IN1(n1886), .IN2(n552), .QN(g10377) );
  INVX0 U1861 ( .IN(n1983), .QN(n1977) );
  INVX0 U1862 ( .IN(n1986), .QN(n1978) );
  INVX0 U1863 ( .IN(n1986), .QN(n1979) );
  INVX0 U1864 ( .IN(n968), .QN(n1952) );
  NAND2X0 U1865 ( .IN1(n797), .IN2(n1395), .QN(n1291) );
  NAND2X0 U1866 ( .IN1(n1974), .IN2(n547), .QN(n1382) );
  INVX0 U1867 ( .IN(n1103), .QN(n557) );
  NAND2X0 U1868 ( .IN1(n668), .IN2(n649), .QN(n1101) );
  NAND2X0 U1869 ( .IN1(n623), .IN2(n715), .QN(n1144) );
  NAND2X0 U1870 ( .IN1(n715), .IN2(n598), .QN(n865) );
  NAND2X0 U1871 ( .IN1(n668), .IN2(n607), .QN(n844) );
  NAND2X0 U1872 ( .IN1(n555), .IN2(n1141), .QN(n1139) );
  NAND2X0 U1873 ( .IN1(n555), .IN2(n661), .QN(n1171) );
  INVX0 U1874 ( .IN(n1984), .QN(n1983) );
  INVX0 U1875 ( .IN(n968), .QN(n1951) );
  INVX0 U1876 ( .IN(n1592), .QN(n592) );
  ISOLANDX1 U1877 ( .D(n1137), .ISO(n1967), .Q(n1195) );
  NOR2X0 U1878 ( .IN1(n1026), .IN2(n649), .QN(n960) );
  NOR2X0 U1879 ( .IN1(n1641), .IN2(n1311), .QN(n1309) );
  INVX0 U1880 ( .IN(n866), .QN(n596) );
  INVX0 U1881 ( .IN(n845), .QN(n606) );
  INVX0 U1882 ( .IN(n850), .QN(n644) );
  INVX0 U1883 ( .IN(n855), .QN(n620) );
  INVX0 U1884 ( .IN(n1407), .QN(n662) );
  NOR2X0 U1885 ( .IN1(n529), .IN2(n1198), .QN(g5763) );
  NOR2X0 U1886 ( .IN1(n533), .IN2(n1181), .QN(g6392) );
  INVX0 U1887 ( .IN(n1005), .QN(n633) );
  INVX0 U1888 ( .IN(n1311), .QN(n611) );
  INVX0 U1889 ( .IN(n1295), .QN(n612) );
  INVX0 U1890 ( .IN(n830), .QN(n603) );
  INVX0 U1891 ( .IN(n875), .QN(n595) );
  INVX0 U1892 ( .IN(n933), .QN(n646) );
  INVX0 U1893 ( .IN(n863), .QN(n712) );
  INVX0 U1894 ( .IN(n908), .QN(n718) );
  AND3X1 U1895 ( .IN1(n1849), .IN2(n1851), .IN3(n1578), .Q(n1575) );
  NAND2X0 U1896 ( .IN1(n1581), .IN2(n1849), .QN(n1579) );
  NAND3X0 U1897 ( .IN1(n1579), .IN2(n1550), .IN3(n1556), .QN(n1473) );
  AND3X1 U1898 ( .IN1(n1831), .IN2(n1841), .IN3(n842), .Q(n1395) );
  AND4X1 U1899 ( .IN1(n1571), .IN2(n583), .IN3(n1572), .IN4(n1573), .Q(n1546)
         );
  NOR2X0 U1900 ( .IN1(n1507), .IN2(n1530), .QN(n1572) );
  NOR4X0 U1901 ( .IN1(n1481), .IN2(n1506), .IN3(n580), .IN4(n1508), .QN(n1573)
         );
  INVX0 U1902 ( .IN(n1239), .QN(n1899) );
  INVX0 U1903 ( .IN(n1900), .QN(n1889) );
  INVX0 U1904 ( .IN(n1239), .QN(n1900) );
  AO21X1 U1905 ( .IN1(n1577), .IN2(n1548), .IN3(n1479), .Q(n1566) );
  XOR3X1 U1906 ( .IN1(n1245), .IN2(n1246), .IN3(n1247), .Q(n1243) );
  XOR2X1 U1907 ( .IN1(n1253), .IN2(n1254), .Q(n1251) );
  ISOLANDX1 U1908 ( .D(n1544), .ISO(n1545), .Q(n1512) );
  ISOLANDX1 U1909 ( .D(n1574), .ISO(n1545), .Q(n1530) );
  AND3X1 U1910 ( .IN1(n1548), .IN2(n1580), .IN3(n1396), .Q(n1859) );
  NAND4X0 U1911 ( .IN1(n1546), .IN2(n1495), .IN3(n1494), .IN4(n1541), .QN(
        n1491) );
  AND2X1 U1912 ( .IN1(n1396), .IN2(n1578), .Q(n1576) );
  XOR2X1 U1913 ( .IN1(n1248), .IN2(n1249), .Q(n1246) );
  NAND4X0 U1914 ( .IN1(n1444), .IN2(n1445), .IN3(n1446), .IN4(n1447), .QN(
        n1440) );
  NAND2X0 U1915 ( .IN1(n1972), .IN2(n1448), .QN(n1446) );
  NAND4X0 U1916 ( .IN1(n547), .IN2(n545), .IN3(n548), .IN4(n1449), .QN(n1448)
         );
  NOR2X0 U1917 ( .IN1(g10663), .IN2(g10664), .QN(n1449) );
  XOR2X1 U1918 ( .IN1(n793), .IN2(n794), .Q(g11163) );
  OA21X1 U1919 ( .IN1(n1302), .IN2(n1606), .IN3(n1903), .Q(n1349) );
  INVX0 U1920 ( .IN(n1239), .QN(n1898) );
  INVX0 U1921 ( .IN(n1239), .QN(n1897) );
  INVX0 U1922 ( .IN(n1239), .QN(n1896) );
  NOR2X0 U1923 ( .IN1(n1344), .IN2(n1345), .QN(g11380) );
  OA21X1 U1924 ( .IN1(n1302), .IN2(n527), .IN3(n1606), .Q(n1344) );
  NOR2X0 U1925 ( .IN1(n1348), .IN2(n1345), .QN(g11372) );
  OA221X1 U1926 ( .IN1(n1349), .IN2(n1594), .IN3(n527), .IN4(n1350), .IN5(
        n1306), .Q(n1348) );
  NAND2X0 U1927 ( .IN1(n1884), .IN2(n1594), .QN(n1350) );
  XOR2X1 U1928 ( .IN1(n544), .IN2(n545), .Q(n1461) );
  XOR3X1 U1929 ( .IN1(n1463), .IN2(n548), .IN3(g10664), .Q(n1462) );
  NOR2X0 U1930 ( .IN1(n1353), .IN2(n1345), .QN(g11340) );
  XOR2X1 U1931 ( .IN1(n527), .IN2(n1884), .Q(n1353) );
  INVX0 U1932 ( .IN(n1464), .QN(g10628) );
  INVX0 U1933 ( .IN(n1541), .QN(n581) );
  NAND4X0 U1934 ( .IN1(n1556), .IN2(n1478), .IN3(n1557), .IN4(n1550), .QN(
        n1552) );
  INVX0 U1935 ( .IN(n1550), .QN(n575) );
  INVX0 U1936 ( .IN(n1495), .QN(n578) );
  INVX0 U1937 ( .IN(n793), .QN(n542) );
  NAND2X0 U1938 ( .IN1(n1974), .IN2(g10664), .QN(n1455) );
  AO221X1 U1939 ( .IN1(n1371), .IN2(g10726), .IN3(n1372), .IN4(g10664), .IN5(
        n1653), .Q(n1369) );
  AO221X1 U1940 ( .IN1(n1373), .IN2(g10720), .IN3(n1374), .IN4(g10722), .IN5(
        n1653), .Q(n1367) );
  AO22X1 U1941 ( .IN1(n662), .IN2(n1069), .IN3(n1454), .IN4(n1407), .Q(n1452)
         );
  NAND2X0 U1942 ( .IN1(n1611), .IN2(n1455), .QN(n1454) );
  AO22X1 U1943 ( .IN1(n662), .IN2(n1075), .IN3(n1404), .IN4(n535), .Q(n1405)
         );
  INVX0 U1944 ( .IN(g10720), .QN(n545) );
  NAND2X0 U1945 ( .IN1(n1973), .IN2(g10721), .QN(n1447) );
  NAND2X0 U1946 ( .IN1(n1968), .IN2(g10719), .QN(n1445) );
  INVX0 U1947 ( .IN(g10724), .QN(n547) );
  INVX0 U1948 ( .IN(g10719), .QN(n544) );
  INVX0 U1949 ( .IN(g10726), .QN(n548) );
  NAND2X0 U1950 ( .IN1(n1969), .IN2(g10720), .QN(n1414) );
  INVX0 U1951 ( .IN(n1987), .QN(n1984) );
  INVX0 U1952 ( .IN(n1987), .QN(n1985) );
  AO22X1 U1953 ( .IN1(n662), .IN2(n1067), .IN3(n1404), .IN4(n532), .Q(n1408)
         );
  AO22X1 U1954 ( .IN1(n662), .IN2(n1063), .IN3(n1418), .IN4(n1407), .Q(n1410)
         );
  NAND2X0 U1955 ( .IN1(n1416), .IN2(n545), .QN(n1418) );
  AO22X1 U1956 ( .IN1(n662), .IN2(n1084), .IN3(n1404), .IN4(n534), .Q(n1412)
         );
  AO22X1 U1957 ( .IN1(n662), .IN2(n1077), .IN3(n1415), .IN4(n1407), .Q(n1411)
         );
  NAND2X0 U1958 ( .IN1(n1416), .IN2(n544), .QN(n1415) );
  INVX0 U1959 ( .IN(g10663), .QN(n552) );
  INVX0 U1960 ( .IN(g10721), .QN(n546) );
  INVX0 U1961 ( .IN(n1255), .QN(n549) );
  AO22X1 U1962 ( .IN1(n662), .IN2(n1082), .IN3(n1413), .IN4(n1407), .Q(n1409)
         );
  NAND2X0 U1963 ( .IN1(n1611), .IN2(n1414), .QN(n1413) );
  XOR2X1 U1964 ( .IN1(g10724), .IN2(g10663), .Q(n1463) );
  NAND2X0 U1965 ( .IN1(n550), .IN2(n1229), .QN(n1225) );
  NAND2X0 U1966 ( .IN1(n1261), .IN2(n1262), .QN(n1259) );
  INVX0 U1967 ( .IN(n1227), .QN(n550) );
  NOR2X0 U1968 ( .IN1(n1965), .IN2(n1113), .QN(n1120) );
  INVX0 U1969 ( .IN(n1867), .QN(n1887) );
  INVX0 U1970 ( .IN(n1867), .QN(n1886) );
  NAND2X0 U1971 ( .IN1(n1113), .IN2(n1114), .QN(n1103) );
  AND4X1 U1972 ( .IN1(n1396), .IN2(n1847), .IN3(n1845), .IN4(n1843), .Q(n797)
         );
  INVX0 U1973 ( .IN(n1988), .QN(n1986) );
  AO221X1 U1974 ( .IN1(n1404), .IN2(g10663), .IN3(n662), .IN4(n1088), .IN5(
        n1450), .Q(n1453) );
  AO22X1 U1975 ( .IN1(n662), .IN2(n1080), .IN3(n1404), .IN4(n1382), .Q(n1402)
         );
  AO221X1 U1976 ( .IN1(n1404), .IN2(g10726), .IN3(n662), .IN4(n1086), .IN5(
        n1450), .Q(n1417) );
  NOR2X0 U1977 ( .IN1(n1217), .IN2(n1961), .QN(g5392) );
  NOR2X0 U1978 ( .IN1(n1683), .IN2(n1961), .QN(n1198) );
  NOR2X0 U1979 ( .IN1(n594), .IN2(n1961), .QN(n1181) );
  NOR2X0 U1980 ( .IN1(n1362), .IN2(n1363), .QN(n1352) );
  NAND2X0 U1981 ( .IN1(n560), .IN2(n744), .QN(n968) );
  INVX0 U1982 ( .IN(n1059), .QN(n533) );
  INVX0 U1983 ( .IN(n1236), .QN(n529) );
  NAND4X0 U1984 ( .IN1(n844), .IN2(n805), .IN3(n952), .IN4(n953), .QN(n845) );
  NOR2X0 U1985 ( .IN1(n954), .IN2(n720), .QN(n952) );
  NAND4X0 U1986 ( .IN1(n865), .IN2(n815), .IN3(n916), .IN4(n715), .QN(n866) );
  ISOLANDX1 U1987 ( .D(n822), .ISO(n809), .Q(n916) );
  NAND4X0 U1988 ( .IN1(n1684), .IN2(n1623), .IN3(n1601), .IN4(n1590), .QN(
        n1289) );
  NAND2X0 U1989 ( .IN1(n648), .IN2(n958), .QN(n850) );
  NAND2X0 U1990 ( .IN1(n622), .IN2(n918), .QN(n855) );
  NAND3X0 U1991 ( .IN1(n1833), .IN2(n1775), .IN3(n842), .QN(g9961) );
  NOR2X0 U1992 ( .IN1(n891), .IN2(n1657), .QN(n875) );
  NOR2X0 U1993 ( .IN1(n949), .IN2(n1656), .QN(n933) );
  NOR2X0 U1994 ( .IN1(n1054), .IN2(n1117), .QN(n1116) );
  NOR2X0 U1995 ( .IN1(n607), .IN2(n805), .QN(n830) );
  NAND2X0 U1996 ( .IN1(n1648), .IN2(n1611), .QN(n1407) );
  NOR2X0 U1997 ( .IN1(n650), .IN2(n954), .QN(n1035) );
  NOR2X0 U1998 ( .IN1(n624), .IN2(n1032), .QN(n1039) );
  NAND2X0 U1999 ( .IN1(n675), .IN2(n1594), .QN(n1311) );
  NAND2X0 U2000 ( .IN1(n985), .IN2(n1658), .QN(n1005) );
  NAND2X0 U2001 ( .IN1(n674), .IN2(n1594), .QN(n1295) );
  NAND2X0 U2002 ( .IN1(n1773), .IN2(n1665), .QN(g8352) );
  NAND2X0 U2003 ( .IN1(n1773), .IN2(n1669), .QN(g8349) );
  NAND2X0 U2004 ( .IN1(n1773), .IN2(n1666), .QN(g8335) );
  NAND2X0 U2005 ( .IN1(n1773), .IN2(n1664), .QN(g8328) );
  NAND2X0 U2006 ( .IN1(n1773), .IN2(n1667), .QN(g8318) );
  NAND2X0 U2007 ( .IN1(n1773), .IN2(n1668), .QN(g8313) );
  NAND2X0 U2008 ( .IN1(n1773), .IN2(n1671), .QN(g8347) );
  NAND2X0 U2009 ( .IN1(n1773), .IN2(n1670), .QN(g8340) );
  NAND2X0 U2010 ( .IN1(n1773), .IN2(n1672), .QN(g8331) );
  NAND2X0 U2011 ( .IN1(n1773), .IN2(n1673), .QN(g8323) );
  NAND2X0 U2012 ( .IN1(n1773), .IN2(n1674), .QN(g8316) );
  NAND3X0 U2013 ( .IN1(n814), .IN2(n815), .IN3(n826), .QN(n863) );
  NAND3X0 U2014 ( .IN1(n831), .IN2(n832), .IN3(n966), .QN(n908) );
  NOR2X0 U2015 ( .IN1(n1029), .IN2(n1622), .QN(n1191) );
  NOR2X0 U2016 ( .IN1(n1593), .IN2(n1607), .QN(n834) );
  NOR2X0 U2017 ( .IN1(n1634), .IN2(n1957), .QN(n1137) );
  INVX0 U2018 ( .IN(n1169), .QN(n538) );
  INVX0 U2019 ( .IN(n1167), .QN(n539) );
  NOR2X0 U2020 ( .IN1(n1963), .IN2(n1159), .QN(n1173) );
  NAND4X0 U2021 ( .IN1(n721), .IN2(n1593), .IN3(n1609), .IN4(n1645), .QN(n1026) );
  NAND4X0 U2022 ( .IN1(n648), .IN2(n718), .IN3(n1615), .IN4(n1662), .QN(n950)
         );
  NAND4X0 U2023 ( .IN1(n622), .IN2(n712), .IN3(n1616), .IN4(n1663), .QN(n892)
         );
  OA221X1 U2024 ( .IN1(n599), .IN2(n810), .IN3(n811), .IN4(n1605), .IN5(n1880), 
        .Q(g9272) );
  NAND2X0 U2025 ( .IN1(n715), .IN2(n1605), .QN(n810) );
  INVX0 U2026 ( .IN(n811), .QN(n599) );
  NAND2X0 U2027 ( .IN1(n812), .IN2(n813), .QN(n811) );
  NOR2X0 U2028 ( .IN1(n1659), .IN2(n1172), .QN(n1141) );
  NOR2X0 U2029 ( .IN1(n1183), .IN2(n1714), .QN(g6179) );
  INVX0 U2030 ( .IN(n1142), .QN(n517) );
  ISOLANDX1 U2031 ( .D(n1057), .ISO(n1054), .Q(n1056) );
  NOR2X0 U2032 ( .IN1(n1626), .IN2(n1117), .QN(n1057) );
  INVX0 U2033 ( .IN(n899), .QN(n648) );
  INVX0 U2034 ( .IN(n853), .QN(n622) );
  ISOLANDX1 U2035 ( .D(n1404), .ISO(n1969), .Q(n1450) );
  OR2X1 U2036 ( .IN1(n1616), .IN2(n922), .Q(n925) );
  OR2X1 U2037 ( .IN1(n1615), .IN2(n846), .Q(n849) );
  NOR2X0 U2038 ( .IN1(n1306), .IN2(n1307), .QN(n1304) );
  NOR3X0 U2039 ( .IN1(n598), .IN2(n1605), .IN3(n826), .QN(n820) );
  NOR2X0 U2040 ( .IN1(n1264), .IN2(n1263), .QN(n1258) );
  AO21X1 U2041 ( .IN1(n605), .IN2(n951), .IN3(n606), .Q(g8883) );
  XOR2X1 U2042 ( .IN1(n1656), .IN2(n955), .Q(n951) );
  NAND2X0 U2043 ( .IN1(n850), .IN2(n956), .QN(n955) );
  NAND3X0 U2044 ( .IN1(n950), .IN2(n949), .IN3(n957), .QN(n956) );
  AO21X1 U2045 ( .IN1(n597), .IN2(n893), .IN3(n596), .Q(g8937) );
  XOR2X1 U2046 ( .IN1(n1657), .IN2(n894), .Q(n893) );
  NAND2X0 U2047 ( .IN1(n855), .IN2(n895), .QN(n894) );
  NAND3X0 U2048 ( .IN1(n892), .IN2(n891), .IN3(n896), .QN(n895) );
  AO21X1 U2049 ( .IN1(n597), .IN2(n887), .IN3(n596), .Q(g8938) );
  XOR2X1 U2050 ( .IN1(n1675), .IN2(n888), .Q(n887) );
  NAND2X0 U2051 ( .IN1(n855), .IN2(n889), .QN(n888) );
  NAND3X0 U2052 ( .IN1(n600), .IN2(n595), .IN3(n890), .QN(n889) );
  AO21X1 U2053 ( .IN1(n605), .IN2(n945), .IN3(n606), .Q(g8885) );
  XOR2X1 U2054 ( .IN1(n1676), .IN2(n946), .Q(n945) );
  NAND2X0 U2055 ( .IN1(n850), .IN2(n947), .QN(n946) );
  NAND3X0 U2056 ( .IN1(n645), .IN2(n646), .IN3(n948), .QN(n947) );
  INVX0 U2057 ( .IN(n1054), .QN(n555) );
  NAND3X0 U2058 ( .IN1(n814), .IN2(n815), .IN3(n816), .QN(n813) );
  OR2X1 U2059 ( .IN1(n817), .IN2(n1643), .Q(n816) );
  NBUFFX2 U2060 ( .IN(n1960), .Q(n1957) );
  NOR2X0 U2061 ( .IN1(n1884), .IN2(n1311), .QN(n1313) );
  NBUFFX2 U2062 ( .IN(n1960), .Q(n1958) );
  NOR2X0 U2063 ( .IN1(n1038), .IN2(n623), .QN(n929) );
  NAND2X0 U2064 ( .IN1(n1593), .IN2(n1644), .QN(n964) );
  NAND2X0 U2065 ( .IN1(n1263), .IN2(n1264), .QN(n1262) );
  NOR2X0 U2066 ( .IN1(n1965), .IN2(n1596), .QN(g4506) );
  NOR2X0 U2067 ( .IN1(n1964), .IN2(n1602), .QN(g6193) );
  NOR2X0 U2068 ( .IN1(n1964), .IN2(n1619), .QN(g6331) );
  NOR2X0 U2069 ( .IN1(n1965), .IN2(n1660), .QN(g4490) );
  NOR2X0 U2070 ( .IN1(n1965), .IN2(n1618), .QN(g4471) );
  NOR2X0 U2071 ( .IN1(n1964), .IN2(n1700), .QN(g6332) );
  NOR2X0 U2072 ( .IN1(n1964), .IN2(n1617), .QN(g4498) );
  NOR2X0 U2073 ( .IN1(n1965), .IN2(n1708), .QN(g4473) );
  NOR2X0 U2074 ( .IN1(n1964), .IN2(n1685), .QN(g4342) );
  NOR2X0 U2075 ( .IN1(n1964), .IN2(n1705), .QN(g4477) );
  NOR2X0 U2076 ( .IN1(n1965), .IN2(n1597), .QN(g4484) );
  NOR2X0 U2077 ( .IN1(n1963), .IN2(n1624), .QN(g6828) );
  NOR2X0 U2078 ( .IN1(n1964), .IN2(n1627), .QN(g6205) );
  NOR2X0 U2079 ( .IN1(n1962), .IN2(n1073), .QN(g8047) );
  XOR2X1 U2080 ( .IN1(n1704), .IN2(g6035), .Q(n1073) );
  NOR2X0 U2081 ( .IN1(n1962), .IN2(n1081), .QN(g8042) );
  XOR2X1 U2082 ( .IN1(n1703), .IN2(n1082), .Q(n1081) );
  NOR2X0 U2083 ( .IN1(n1963), .IN2(n1625), .QN(g6820) );
  NOR2X0 U2084 ( .IN1(n1963), .IN2(n1603), .QN(g6334) );
  NOR2X0 U2085 ( .IN1(n1965), .IN2(n1661), .QN(g4465) );
  NOR2X0 U2086 ( .IN1(n1963), .IN2(n1688), .QN(g6834) );
  NOR2X0 U2087 ( .IN1(n1963), .IN2(n1598), .QN(g6840) );
  NOR2X0 U2088 ( .IN1(n1964), .IN2(n1628), .QN(g6180) );
  NOR2X0 U2089 ( .IN1(n1965), .IN2(n1706), .QN(g4480) );
  NOR2X0 U2090 ( .IN1(n1964), .IN2(n1710), .QN(g6224) );
  NOR2X0 U2091 ( .IN1(n1963), .IN2(n1711), .QN(g6839) );
  NOR2X0 U2092 ( .IN1(n1964), .IN2(n1678), .QN(g6333) );
  NOR2X0 U2093 ( .IN1(n1963), .IN2(n1629), .QN(g6841) );
  NOR2X0 U2094 ( .IN1(n1965), .IN2(n1686), .QN(g4340) );
  NOR2X0 U2095 ( .IN1(n1963), .IN2(n1687), .QN(g6830) );
  NOR2X0 U2096 ( .IN1(n1953), .IN2(n1648), .QN(g4500) );
  NOR2X0 U2097 ( .IN1(n1654), .IN2(n1216), .QN(g5390) );
  NOR2X0 U2098 ( .IN1(n1614), .IN2(n1216), .QN(g5148) );
  NOR2X0 U2099 ( .IN1(n1677), .IN2(n1216), .QN(g5173) );
  NOR2X0 U2100 ( .IN1(n1658), .IN2(n1216), .QN(g5126) );
  NOR2X0 U2101 ( .IN1(n1630), .IN2(n1040), .QN(g8254) );
  NOR2X0 U2102 ( .IN1(n1604), .IN2(n1040), .QN(g8147) );
  NOR2X0 U2103 ( .IN1(n1591), .IN2(n1040), .QN(g8250) );
  NOR2X0 U2104 ( .IN1(n1712), .IN2(n1040), .QN(g8260) );
  NOR2X0 U2105 ( .IN1(n644), .IN2(n912), .QN(n911) );
  NOR2X0 U2106 ( .IN1(n620), .IN2(n869), .QN(n868) );
  NBUFFX2 U2107 ( .IN(n1960), .Q(n1959) );
  NAND2X0 U2108 ( .IN1(n830), .IN2(n1713), .QN(n803) );
  NAND2X0 U2109 ( .IN1(n685), .IN2(n1595), .QN(n1128) );
  INVX0 U2110 ( .IN(n1183), .QN(n519) );
  NOR3X0 U2111 ( .IN1(n1953), .IN2(g4089), .IN3(n561), .QN(g5083) );
  NOR2X0 U2112 ( .IN1(n1885), .IN2(n1170), .QN(g6516) );
  OA22X1 U2113 ( .IN1(n1141), .IN2(n1171), .IN3(n554), .IN4(n1659), .Q(n1170)
         );
  INVX0 U2114 ( .IN(n1139), .QN(n554) );
  NOR2X0 U2115 ( .IN1(n1885), .IN2(n1115), .QN(g7541) );
  OA22X1 U2116 ( .IN1(n1057), .IN2(n556), .IN3(n1056), .IN4(n1626), .Q(n1115)
         );
  INVX0 U2117 ( .IN(n1116), .QN(n556) );
  NAND2X0 U2118 ( .IN1(n1605), .IN2(n1643), .QN(n928) );
  NOR2X0 U2119 ( .IN1(n1957), .IN2(n839), .QN(g9110) );
  XOR2X1 U2120 ( .IN1(n1607), .IN2(n840), .Q(n839) );
  NAND3X0 U2121 ( .IN1(n837), .IN2(n603), .IN3(n841), .QN(n840) );
  NAND2X0 U2122 ( .IN1(n804), .IN2(n719), .QN(n841) );
  INVX0 U2123 ( .IN(n1160), .QN(n667) );
  INVX0 U2124 ( .IN(n1148), .QN(n711) );
  NAND2X0 U2125 ( .IN1(n1160), .IN2(n1701), .QN(g6672) );
  NAND2X0 U2126 ( .IN1(n795), .IN2(n796), .QN(n1585) );
  NAND2X0 U2127 ( .IN1(n797), .IN2(n798), .QN(n1587) );
  NAND2X0 U2128 ( .IN1(n795), .IN2(n798), .QN(n1588) );
  NAND2X0 U2129 ( .IN1(n797), .IN2(n796), .QN(n1586) );
  INVX0 U2130 ( .IN(n1016), .QN(n650) );
  INVX0 U2131 ( .IN(n1031), .QN(n624) );
  NAND4X0 U2132 ( .IN1(n1380), .IN2(n822), .IN3(n1038), .IN4(n920), .QN(n1379)
         );
  NAND2X0 U2133 ( .IN1(n713), .IN2(n1605), .QN(n814) );
  NAND2X0 U2134 ( .IN1(n719), .IN2(n1593), .QN(n831) );
  INVX0 U2135 ( .IN(n1046), .QN(n537) );
  INVX0 U2136 ( .IN(n1025), .QN(n719) );
  INVX0 U2137 ( .IN(n1306), .QN(n610) );
  INVX0 U2138 ( .IN(n978), .QN(n631) );
  INVX0 U2139 ( .IN(n954), .QN(n668) );
  INVX0 U2140 ( .IN(n1109), .QN(n540) );
  INVX0 U2141 ( .IN(n1032), .QN(n715) );
  INVX0 U2142 ( .IN(n1325), .QN(n674) );
  INVX0 U2143 ( .IN(n1307), .QN(n675) );
  INVX0 U2144 ( .IN(n920), .QN(n713) );
  INVX0 U2145 ( .IN(n877), .QN(n600) );
  INVX0 U2146 ( .IN(n935), .QN(n645) );
  INVX0 U2147 ( .IN(n1092), .QN(n630) );
  INVX0 U2148 ( .IN(n953), .QN(n717) );
  OAI21X1 U2149 ( .IN1(n915), .IN2(n865), .IN3(n866), .QN(g8921) );
  OA22X1 U2150 ( .IN1(n922), .IN2(n923), .IN3(n924), .IN4(n1616), .Q(n915) );
  NAND2X0 U2151 ( .IN1(n855), .IN2(n925), .QN(n923) );
  NOR2X0 U2152 ( .IN1(n620), .IN2(n925), .QN(n924) );
  OAI21X1 U2153 ( .IN1(n843), .IN2(n844), .IN3(n845), .QN(g8973) );
  OA22X1 U2154 ( .IN1(n846), .IN2(n847), .IN3(n848), .IN4(n1615), .Q(n843) );
  NAND2X0 U2155 ( .IN1(n850), .IN2(n849), .QN(n847) );
  NOR2X0 U2156 ( .IN1(n644), .IN2(n849), .QN(n848) );
  OAI21X1 U2157 ( .IN1(n909), .IN2(n844), .IN3(n845), .QN(g8922) );
  OA22X1 U2158 ( .IN1(n647), .IN2(n910), .IN3(n911), .IN4(n1662), .Q(n909) );
  INVX0 U2159 ( .IN(n913), .QN(n647) );
  NAND2X0 U2160 ( .IN1(n850), .IN2(n912), .QN(n910) );
  OAI21X1 U2161 ( .IN1(n864), .IN2(n865), .IN3(n866), .QN(g8943) );
  OA22X1 U2162 ( .IN1(n621), .IN2(n867), .IN3(n868), .IN4(n1663), .Q(n864) );
  INVX0 U2163 ( .IN(n870), .QN(n621) );
  NAND2X0 U2164 ( .IN1(n855), .IN2(n869), .QN(n867) );
  INVX0 U2165 ( .IN(n1384), .QN(n536) );
  INVX0 U2166 ( .IN(n1042), .QN(n520) );
  INVX0 U2167 ( .IN(n1119), .QN(n685) );
  OA221X1 U2168 ( .IN1(n604), .IN2(n827), .IN3(n828), .IN4(n1593), .IN5(g2355), 
        .Q(g9150) );
  NAND2X0 U2169 ( .IN1(n668), .IN2(n1593), .QN(n827) );
  INVX0 U2170 ( .IN(n828), .QN(n604) );
  OA21X1 U2171 ( .IN1(n607), .IN2(n829), .IN3(n803), .Q(n828) );
  INVX0 U2172 ( .IN(n966), .QN(n721) );
  INVX0 U2173 ( .IN(n959), .QN(n649) );
  INVX0 U2174 ( .IN(n993), .QN(n632) );
  INVX0 U2175 ( .IN(n1318), .QN(n609) );
  INVX0 U2176 ( .IN(n999), .QN(n634) );
  INVX0 U2177 ( .IN(n926), .QN(n623) );
  INVX0 U2178 ( .IN(n832), .QN(n720) );
  INVX0 U2179 ( .IN(n1302), .QN(n614) );
  INVX0 U2180 ( .IN(n804), .QN(n607) );
  INVX0 U2181 ( .IN(n812), .QN(n598) );
  INVX0 U2182 ( .IN(n1114), .QN(n629) );
  INVX0 U2183 ( .IN(n1110), .QN(n665) );
  INVX0 U2184 ( .IN(n974), .QN(n564) );
  INVX0 U2185 ( .IN(n995), .QN(n568) );
  INVX0 U2186 ( .IN(n1001), .QN(n566) );
  INVX0 U2187 ( .IN(n981), .QN(n563) );
  INVX0 U2188 ( .IN(n989), .QN(n567) );
  INVX0 U2189 ( .IN(n1007), .QN(n569) );
  INVX0 U2190 ( .IN(n1012), .QN(n565) );
  INVX0 U2191 ( .IN(n1420), .QN(n625) );
  INVX0 U2192 ( .IN(n1166), .QN(n518) );
  INVX0 U2193 ( .IN(n1875), .QN(n1888) );
  NOR2X0 U2194 ( .IN1(n1126), .IN2(n1101), .QN(g7137) );
  OA22X1 U2195 ( .IN1(n1127), .IN2(n1709), .IN3(n651), .IN4(n1128), .Q(n1126)
         );
  INVX0 U2196 ( .IN(n1129), .QN(n651) );
  NOR2X0 U2197 ( .IN1(n1701), .IN2(n1129), .QN(n1127) );
  NOR2X0 U2198 ( .IN1(n1130), .IN2(n1101), .QN(g7134) );
  OA21X1 U2199 ( .IN1(n685), .IN2(n1595), .IN3(n1128), .Q(n1130) );
  INVX0 U2200 ( .IN(n1217), .QN(n725) );
  NOR4X0 U2201 ( .IN1(n1712), .IN2(n1630), .IN3(n1604), .IN4(n1591), .QN(g3381) );
  NOR2X0 U2202 ( .IN1(n592), .IN2(n1664), .QN(g6638) );
  NOR2X0 U2203 ( .IN1(n592), .IN2(n1665), .QN(g6531) );
  NOR2X0 U2204 ( .IN1(n592), .IN2(n1666), .QN(g6653) );
  NOR2X0 U2205 ( .IN1(n592), .IN2(n1667), .QN(g6627) );
  NOR2X0 U2206 ( .IN1(n592), .IN2(n1668), .QN(g6621) );
  NOR2X0 U2207 ( .IN1(n592), .IN2(n1669), .QN(g6526) );
  NAND2X0 U2208 ( .IN1(n1148), .IN2(n1642), .QN(g6755) );
  NOR2X0 U2209 ( .IN1(n555), .IN2(n1601), .QN(g10780) );
  NOR2X0 U2210 ( .IN1(n555), .IN2(n1623), .QN(g10785) );
  NOR2X0 U2211 ( .IN1(n555), .IN2(n1684), .QN(g10784) );
  NOR2X0 U2212 ( .IN1(n555), .IN2(n1590), .QN(g10782) );
  INVX0 U2213 ( .IN(n1451), .QN(n561) );
  NAND2X0 U2214 ( .IN1(n1670), .IN2(n1592), .QN(g7219) );
  NAND2X0 U2215 ( .IN1(n1671), .IN2(n1592), .QN(g7143) );
  NAND2X0 U2216 ( .IN1(n1672), .IN2(n1592), .QN(g7204) );
  NAND2X0 U2217 ( .IN1(n1673), .IN2(n1592), .QN(g7189) );
  NAND2X0 U2218 ( .IN1(n1674), .IN2(n1592), .QN(g7183) );
  INVX0 U2219 ( .IN(n1228), .QN(n687) );
  INVX0 U2220 ( .IN(n1338), .QN(n616) );
  INVX0 U2221 ( .IN(n1342), .QN(n617) );
  INVX0 U2222 ( .IN(n1172), .QN(n661) );
  OA22X1 U2223 ( .IN1(n577), .IN2(n1632), .IN3(n583), .IN4(DFF_228_n1), .Q(
        n1499) );
  AOI221X1 U2224 ( .IN1(n1479), .IN2(g1558), .IN3(n1480), .IN4(g1601), .IN5(
        n1513), .QN(n1501) );
  NAND2X0 U2225 ( .IN1(g6257), .IN2(n1581), .QN(n1550) );
  NOR3X0 U2226 ( .IN1(g833), .IN2(g841), .IN3(g837), .QN(n1441) );
  NOR4X0 U2227 ( .IN1(n1443), .IN2(g853), .IN3(g861), .IN4(g857), .QN(n1442)
         );
  NAND2X0 U2228 ( .IN1(g6263), .IN2(n1775), .QN(n1484) );
  NAND2X0 U2229 ( .IN1(n1547), .IN2(g6257), .QN(n1495) );
  NOR2X0 U2230 ( .IN1(n1849), .IN2(g6258), .QN(n1396) );
  NOR2X0 U2231 ( .IN1(g6263), .IN2(g6256), .QN(n1583) );
  NOR2X0 U2232 ( .IN1(n1847), .IN2(g6260), .QN(n1580) );
  AND4X1 U2233 ( .IN1(n1548), .IN2(g6258), .IN3(n1847), .IN4(n1845), .Q(n1547)
         );
  AND3X1 U2234 ( .IN1(n842), .IN2(n1831), .IN3(g6262), .Q(n796) );
  AND3X1 U2235 ( .IN1(n842), .IN2(n1841), .IN3(g6261), .Q(n798) );
  NOR2X0 U2236 ( .IN1(n1845), .IN2(g6259), .QN(n1578) );
  NOR2X0 U2237 ( .IN1(n1843), .IN2(g6256), .QN(n1569) );
  AND3X1 U2238 ( .IN1(g6257), .IN2(g6258), .IN3(n1580), .Q(n1577) );
  AO222X1 U2239 ( .IN1(n572), .IN2(g1753), .IN3(n579), .IN4(n1631), .IN5(n575), 
        .IN6(g1730), .Q(n1513) );
  AO21X1 U2240 ( .IN1(g318), .IN2(n1905), .IN3(n1315), .Q(n1247) );
  OA221X1 U2241 ( .IN1(n1316), .IN2(g486), .IN3(n1621), .IN4(n1317), .IN5(
        n1902), .Q(n1315) );
  NAND2X0 U2242 ( .IN1(n609), .IN2(n1883), .QN(n1317) );
  NOR2X0 U2243 ( .IN1(n1641), .IN2(n1318), .QN(n1316) );
  AO21X1 U2244 ( .IN1(g330), .IN2(n1904), .IN3(n1299), .Q(n1252) );
  OA221X1 U2245 ( .IN1(n1300), .IN2(g506), .IN3(n1600), .IN4(n1301), .IN5(
        n1854), .Q(n1299) );
  NAND2X0 U2246 ( .IN1(n614), .IN2(n1606), .QN(n1301) );
  NOR2X0 U2247 ( .IN1(g471), .IN2(n1302), .QN(n1300) );
  AO22X1 U2248 ( .IN1(n1592), .IN2(g336), .IN3(n1219), .IN4(n592), .Q(g11647)
         );
  OAI22X1 U2249 ( .IN1(n551), .IN2(n1220), .IN3(n1221), .IN4(n1222), .QN(n1219) );
  INVX0 U2250 ( .IN(n1222), .QN(n551) );
  AO22X1 U2251 ( .IN1(g345), .IN2(n1592), .IN3(n1237), .IN4(n592), .Q(g11625)
         );
  XOR2X1 U2252 ( .IN1(n1220), .IN2(n1221), .Q(n1237) );
  AO21X1 U2253 ( .IN1(g324), .IN2(n1906), .IN3(n1308), .Q(n1249) );
  OA221X1 U2254 ( .IN1(n1309), .IN2(g496), .IN3(n1689), .IN4(n1310), .IN5(
        n1901), .Q(n1308) );
  NAND2X0 U2255 ( .IN1(n611), .IN2(n1884), .QN(n1310) );
  AO21X1 U2256 ( .IN1(g309), .IN2(n1904), .IN3(n1292), .Q(n1254) );
  OA221X1 U2257 ( .IN1(n1293), .IN2(g516), .IN3(n1620), .IN4(n1294), .IN5(
        n1901), .Q(n1292) );
  NAND2X0 U2258 ( .IN1(n1884), .IN2(n612), .QN(n1294) );
  NOR2X0 U2259 ( .IN1(n1295), .IN2(n1641), .QN(n1293) );
  AO21X1 U2260 ( .IN1(g315), .IN2(n1907), .IN3(n1319), .Q(n1245) );
  OA221X1 U2261 ( .IN1(n1320), .IN2(g481), .IN3(n1680), .IN4(n1321), .IN5(
        n1901), .Q(n1319) );
  NAND2X0 U2262 ( .IN1(n609), .IN2(n1641), .QN(n1321) );
  NOR2X0 U2263 ( .IN1(n1884), .IN2(n1318), .QN(n1320) );
  AO21X1 U2264 ( .IN1(g327), .IN2(n1905), .IN3(n1303), .Q(n1250) );
  OA221X1 U2265 ( .IN1(n1304), .IN2(g501), .IN3(n1690), .IN4(n1305), .IN5(
        n1901), .Q(n1303) );
  NAND2X0 U2266 ( .IN1(n675), .IN2(n610), .QN(n1305) );
  AO21X1 U2267 ( .IN1(g321), .IN2(n1908), .IN3(n1312), .Q(n1248) );
  OA221X1 U2268 ( .IN1(n1313), .IN2(g491), .IN3(n1691), .IN4(n1314), .IN5(
        n1901), .Q(n1312) );
  NAND2X0 U2269 ( .IN1(n611), .IN2(n1641), .QN(n1314) );
  AO21X1 U2270 ( .IN1(g333), .IN2(n1906), .IN3(n1296), .Q(n1253) );
  OA221X1 U2271 ( .IN1(n1297), .IN2(g511), .IN3(n1679), .IN4(n1298), .IN5(
        n1901), .Q(n1296) );
  NAND2X0 U2272 ( .IN1(n612), .IN2(n1641), .QN(n1298) );
  NOR2X0 U2273 ( .IN1(n1884), .IN2(n1295), .QN(n1297) );
  NOR3X0 U2274 ( .IN1(n1503), .IN2(n1504), .IN3(n1505), .QN(n1502) );
  AO222X1 U2275 ( .IN1(g986), .IN2(n1506), .IN3(g959), .IN4(n580), .IN5(g4199), 
        .IN6(n1481), .Q(n1505) );
  AOI22X1 U2276 ( .IN1(n1506), .IN2(g947), .IN3(n1483), .IN4(g284), .QN(n1553)
         );
  OA221X1 U2277 ( .IN1(n583), .IN2(DFF_319_n1), .IN3(n1550), .IN4(n1633), 
        .IN5(n1555), .Q(n1554) );
  NOR2X0 U2278 ( .IN1(n1545), .IN2(n1831), .QN(n1570) );
  AOI22X1 U2279 ( .IN1(n1860), .IN2(n1861), .IN3(n1861), .IN4(n1459), .QN(n793) );
  OR2X1 U2280 ( .IN1(g32), .IN2(n583), .Q(n1860) );
  OAI21X1 U2281 ( .IN1(g32), .IN2(n583), .IN3(n1459), .QN(n1861) );
  AO221X1 U2282 ( .IN1(g5392), .IN2(g10663), .IN3(n535), .IN4(n1198), .IN5(
        n1465), .Q(n794) );
  AO222X1 U2283 ( .IN1(n1466), .IN2(n1977), .IN3(g2648), .IN4(n530), .IN5(n529), .IN6(g10724), .Q(n1465) );
  NOR2X0 U2284 ( .IN1(g105), .IN2(n548), .QN(n1466) );
  INVX0 U2285 ( .IN(n1455), .QN(n530) );
  NAND3X0 U2286 ( .IN1(n1853), .IN2(n1419), .IN3(n1420), .QN(n1337) );
  NAND4X0 U2287 ( .IN1(n1421), .IN2(n1422), .IN3(n1423), .IN4(n1424), .QN(
        n1419) );
  XNOR2X1 U2288 ( .IN1(g330), .IN2(g406), .Q(n1421) );
  XNOR2X1 U2289 ( .IN1(g309), .IN2(g416), .Q(n1422) );
  AO22X1 U2290 ( .IN1(g305), .IN2(n1910), .IN3(n1238), .IN4(n1903), .Q(n1221)
         );
  XNOR2X1 U2291 ( .IN1(n1240), .IN2(n1241), .Q(n1238) );
  NAND4X0 U2292 ( .IN1(n1884), .IN2(n1594), .IN3(n1646), .IN4(n1606), .QN(
        n1240) );
  AO221X1 U2293 ( .IN1(n1181), .IN2(g10720), .IN3(n1362), .IN4(g10724), .IN5(
        n1467), .Q(n1464) );
  AO222X1 U2294 ( .IN1(n1363), .IN2(n535), .IN3(g877), .IN4(n534), .IN5(n533), 
        .IN6(n532), .Q(n1467) );
  AO22X1 U2295 ( .IN1(g516), .IN2(n1902), .IN3(n1911), .IN4(g476), .Q(g11338)
         );
  AO22X1 U2296 ( .IN1(g506), .IN2(n1854), .IN3(g511), .IN4(n1911), .Q(g11336)
         );
  AO22X1 U2297 ( .IN1(g538), .IN2(n1854), .IN3(g534), .IN4(n1911), .Q(g11327)
         );
  AO22X1 U2298 ( .IN1(g530), .IN2(n1853), .IN3(g525), .IN4(n1913), .Q(g11329)
         );
  AO22X1 U2299 ( .IN1(g501), .IN2(n1902), .IN3(g506), .IN4(n1915), .Q(g11335)
         );
  AO22X1 U2300 ( .IN1(g525), .IN2(n1854), .IN3(g521), .IN4(n1913), .Q(g11330)
         );
  AO22X1 U2301 ( .IN1(n1241), .IN2(n1853), .IN3(g481), .IN4(n1914), .Q(g11324)
         );
  AO22X1 U2302 ( .IN1(g416), .IN2(n1902), .IN3(g421), .IN4(n1918), .Q(g11270)
         );
  AO22X1 U2303 ( .IN1(g486), .IN2(n1854), .IN3(g491), .IN4(n1912), .Q(g11332)
         );
  AO22X1 U2304 ( .IN1(g511), .IN2(n1853), .IN3(g516), .IN4(n1911), .Q(g11337)
         );
  AO22X1 U2305 ( .IN1(g496), .IN2(n1902), .IN3(g501), .IN4(n1912), .Q(g11334)
         );
  AO22X1 U2306 ( .IN1(g534), .IN2(n1853), .IN3(g530), .IN4(n1911), .Q(g11328)
         );
  AO22X1 U2307 ( .IN1(g476), .IN2(n1902), .IN3(g542), .IN4(n1915), .Q(g11325)
         );
  AO22X1 U2308 ( .IN1(g411), .IN2(n1854), .IN3(g416), .IN4(n1917), .Q(g11269)
         );
  AO22X1 U2309 ( .IN1(g542), .IN2(n1853), .IN3(g538), .IN4(n1916), .Q(g11326)
         );
  AO22X1 U2310 ( .IN1(g481), .IN2(n1902), .IN3(g486), .IN4(n1912), .Q(g11331)
         );
  AO22X1 U2311 ( .IN1(g391), .IN2(n1854), .IN3(g396), .IN4(n1918), .Q(g11265)
         );
  AO22X1 U2312 ( .IN1(g491), .IN2(n1853), .IN3(g496), .IN4(n1916), .Q(g11333)
         );
  AO22X1 U2313 ( .IN1(g440), .IN2(n1903), .IN3(g435), .IN4(n1920), .Q(g11261)
         );
  AO22X1 U2314 ( .IN1(g435), .IN2(n1903), .IN3(g431), .IN4(n1921), .Q(g11262)
         );
  AO22X1 U2315 ( .IN1(g406), .IN2(n1903), .IN3(g411), .IN4(n1917), .Q(g11268)
         );
  AO22X1 U2316 ( .IN1(g401), .IN2(n1903), .IN3(g406), .IN4(n1916), .Q(g11267)
         );
  AO22X1 U2317 ( .IN1(g386), .IN2(n1903), .IN3(g391), .IN4(n1918), .Q(g11264)
         );
  AO22X1 U2318 ( .IN1(g444), .IN2(n1903), .IN3(g440), .IN4(n1920), .Q(g11260)
         );
  AO22X1 U2319 ( .IN1(g452), .IN2(n1903), .IN3(g448), .IN4(n1910), .Q(g11258)
         );
  AO22X1 U2320 ( .IN1(g426), .IN2(n1903), .IN3(g386), .IN4(n1918), .Q(g11263)
         );
  AO22X1 U2321 ( .IN1(g396), .IN2(n1903), .IN3(g401), .IN4(n1919), .Q(g11266)
         );
  AO22X1 U2322 ( .IN1(g448), .IN2(n1903), .IN3(g444), .IN4(n1919), .Q(g11259)
         );
  AO22X1 U2323 ( .IN1(n602), .IN2(n1903), .IN3(g426), .IN4(n1914), .Q(g11256)
         );
  INVX0 U2324 ( .IN(n1390), .QN(n602) );
  AO22X1 U2325 ( .IN1(g421), .IN2(n1903), .IN3(g452), .IN4(n1921), .Q(g11257)
         );
  AO22X1 U2326 ( .IN1(g833), .IN2(n1855), .IN3(g947), .IN4(n1361), .Q(g11300)
         );
  AO22X1 U2327 ( .IN1(g845), .IN2(n1855), .IN3(g956), .IN4(n1361), .Q(g11306)
         );
  AO22X1 U2328 ( .IN1(g837), .IN2(n1855), .IN3(g950), .IN4(n1361), .Q(g11303)
         );
  AO22X1 U2329 ( .IN1(g861), .IN2(n1855), .IN3(g968), .IN4(n1361), .Q(g11314)
         );
  AO22X1 U2330 ( .IN1(g841), .IN2(n1855), .IN3(g953), .IN4(n1361), .Q(g11305)
         );
  AO22X1 U2331 ( .IN1(g829), .IN2(n1855), .IN3(g944), .IN4(n1361), .Q(g11298)
         );
  AO22X1 U2332 ( .IN1(g857), .IN2(n1855), .IN3(g965), .IN4(n1361), .Q(g11312)
         );
  AO22X1 U2333 ( .IN1(g853), .IN2(n1855), .IN3(g962), .IN4(n1361), .Q(g11310)
         );
  AO22X1 U2334 ( .IN1(g849), .IN2(n1855), .IN3(g959), .IN4(n1361), .Q(g11308)
         );
  AO22X1 U2335 ( .IN1(g339), .IN2(n1592), .IN3(n592), .IN4(n1244), .Q(g11478)
         );
  AO22X1 U2336 ( .IN1(g363), .IN2(n1592), .IN3(n592), .IN4(n1252), .Q(g11486)
         );
  AO22X1 U2337 ( .IN1(g351), .IN2(n1592), .IN3(n592), .IN4(n1247), .Q(g11482)
         );
  AO22X1 U2338 ( .IN1(g348), .IN2(n1592), .IN3(n592), .IN4(n1245), .Q(g11481)
         );
  AO22X1 U2339 ( .IN1(g366), .IN2(n1592), .IN3(n592), .IN4(n1253), .Q(g11487)
         );
  AO22X1 U2340 ( .IN1(g360), .IN2(n1592), .IN3(n592), .IN4(n1250), .Q(g11485)
         );
  AO22X1 U2341 ( .IN1(g342), .IN2(n1592), .IN3(n592), .IN4(n1254), .Q(g11488)
         );
  AO22X1 U2342 ( .IN1(g357), .IN2(n1592), .IN3(n592), .IN4(n1249), .Q(g11484)
         );
  AO22X1 U2343 ( .IN1(g354), .IN2(n1592), .IN3(n592), .IN4(n1248), .Q(g11483)
         );
  AO21X1 U2344 ( .IN1(g312), .IN2(n1907), .IN3(n1322), .Q(n1244) );
  OA221X1 U2345 ( .IN1(n1323), .IN2(g476), .IN3(n1599), .IN4(n1324), .IN5(
        n1854), .Q(n1322) );
  NAND2X0 U2346 ( .IN1(n610), .IN2(n674), .QN(n1324) );
  NOR2X0 U2347 ( .IN1(n1325), .IN2(n1306), .QN(n1323) );
  NOR2X0 U2348 ( .IN1(n1333), .IN2(n1334), .QN(g11393) );
  OA22X1 U2349 ( .IN1(n616), .IN2(n1335), .IN3(n1336), .IN4(n1722), .Q(n1333)
         );
  NOR2X0 U2350 ( .IN1(n1337), .IN2(n1338), .QN(n1336) );
  NOR2X0 U2351 ( .IN1(n1339), .IN2(n1334), .QN(g11392) );
  OA22X1 U2352 ( .IN1(n1340), .IN2(n1341), .IN3(n522), .IN4(n1720), .Q(n1339)
         );
  NAND2X0 U2353 ( .IN1(g976), .IN2(n1342), .QN(n1341) );
  NOR2X0 U2354 ( .IN1(n1343), .IN2(n1334), .QN(g11391) );
  XOR2X1 U2355 ( .IN1(n1340), .IN2(g976), .Q(n1343) );
  NOR2X0 U2356 ( .IN1(n1359), .IN2(n536), .QN(g11320) );
  XOR2X1 U2357 ( .IN1(g369), .IN2(n1360), .Q(n1359) );
  NOR2X0 U2358 ( .IN1(n1351), .IN2(n1334), .QN(g11349) );
  XOR2X1 U2359 ( .IN1(g971), .IN2(n1337), .Q(n1351) );
  OA21X1 U2360 ( .IN1(n1346), .IN2(n1347), .IN3(n521), .Q(g11376) );
  INVX0 U2361 ( .IN(n1345), .QN(n521) );
  OA21X1 U2362 ( .IN1(n1302), .IN2(n527), .IN3(g466), .Q(n1347) );
  NOR4X0 U2363 ( .IN1(n614), .IN2(n1594), .IN3(n1641), .IN4(n527), .QN(n1346)
         );
  OA21X1 U2364 ( .IN1(n1383), .IN2(g382), .IN3(n1384), .Q(g11292) );
  NOR2X0 U2365 ( .IN1(n1385), .IN2(n1360), .QN(n1383) );
  OA21X1 U2366 ( .IN1(n1386), .IN2(n1387), .IN3(n1384), .Q(g11291) );
  OA21X1 U2367 ( .IN1(n1385), .IN2(n1360), .IN3(g378), .Q(n1387) );
  AND4X1 U2368 ( .IN1(n1385), .IN2(g369), .IN3(g374), .IN4(n526), .Q(n1386) );
  NAND2X0 U2369 ( .IN1(n524), .IN2(g971), .QN(n1340) );
  NOR2X0 U2370 ( .IN1(n1388), .IN2(n536), .QN(g11290) );
  XOR2X1 U2371 ( .IN1(n1389), .IN2(g374), .Q(n1388) );
  AO22X1 U2372 ( .IN1(g1669), .IN2(n1888), .IN3(n1403), .IN4(n1404), .Q(g10865) );
  OA21X1 U2373 ( .IN1(g10722), .IN2(n1966), .IN3(n1875), .Q(n1403) );
  AO22X1 U2374 ( .IN1(n561), .IN2(n535), .IN3(g1730), .IN4(n1451), .Q(g10707)
         );
  AO22X1 U2375 ( .IN1(n1875), .IN2(n1452), .IN3(g1657), .IN4(n1888), .Q(g10767) );
  AO22X1 U2376 ( .IN1(g560), .IN2(n1930), .IN3(n1954), .IN4(n1405), .Q(g10797)
         );
  AO22X1 U2377 ( .IN1(g1681), .IN2(n1929), .IN3(n1955), .IN4(n1405), .Q(g10864) );
  AO22X1 U2378 ( .IN1(g572), .IN2(n1930), .IN3(n1954), .IN4(n1452), .Q(g10718)
         );
  AO221X1 U2379 ( .IN1(n1032), .IN2(n1364), .IN3(n619), .IN4(g1857), .IN5(
        n1365), .Q(g11294) );
  AND3X1 U2380 ( .IN1(n1366), .IN2(n1682), .IN3(n926), .Q(n1365) );
  NAND4X0 U2381 ( .IN1(n1367), .IN2(n1368), .IN3(n1369), .IN4(n1370), .QN(
        n1364) );
  NAND4X0 U2382 ( .IN1(n815), .IN2(n822), .IN3(n920), .IN4(n817), .QN(n1366)
         );
  AO22X1 U2383 ( .IN1(g1811), .IN2(n1054), .IN3(n555), .IN4(n1391), .Q(g10936)
         );
  NAND4X0 U2384 ( .IN1(n1291), .IN2(n547), .IN3(n535), .IN4(n1392), .QN(n1391)
         );
  AND3X1 U2385 ( .IN1(n545), .IN2(n544), .IN3(n546), .Q(n1392) );
  NAND4X0 U2386 ( .IN1(n1523), .IN2(n1524), .IN3(n1525), .IN4(n1526), .QN(
        g10720) );
  AOI222X1 U2387 ( .IN1(n1479), .IN2(g1552), .IN3(n572), .IN4(g1747), .IN5(
        n1480), .IN6(g1595), .QN(n1523) );
  AOI222X1 U2388 ( .IN1(n575), .IN2(g1724), .IN3(n578), .IN4(g4), .IN5(n579), 
        .IN6(g12), .QN(n1524) );
  OA221X1 U2389 ( .IN1(n583), .IN2(DFF_384_n1), .IN3(n577), .IN4(n1635), .IN5(
        n1532), .Q(n1525) );
  NOR3X0 U2390 ( .IN1(n1527), .IN2(n1528), .IN3(n1529), .QN(n1526) );
  AO222X1 U2391 ( .IN1(g953), .IN2(n580), .IN3(g932), .IN4(n1508), .IN5(g976), 
        .IN6(n1506), .Q(n1529) );
  NAND4X0 U2392 ( .IN1(n1558), .IN2(n1559), .IN3(n1560), .IN4(n1561), .QN(
        g10663) );
  NOR4X0 U2393 ( .IN1(n1562), .IN2(n1563), .IN3(n581), .IN4(n1564), .QN(n1561)
         );
  AOI22X1 U2394 ( .IN1(n572), .IN2(g1762), .IN3(n1483), .IN4(g281), .QN(n1558)
         );
  AOI222X1 U2395 ( .IN1(n1484), .IN2(n1637), .IN3(n1485), .IN4(g1586), .IN5(
        n1486), .IN6(g1543), .QN(n1560) );
  NAND4X0 U2396 ( .IN1(n1487), .IN2(n1488), .IN3(n1489), .IN4(n1490), .QN(
        g10724) );
  OA221X1 U2397 ( .IN1(n1494), .IN2(DFF_122_n1), .IN3(n1495), .IN4(DFF_445_n1), 
        .IN5(n1496), .Q(n1489) );
  AOI221X1 U2398 ( .IN1(n1483), .IN2(g275), .IN3(n1482), .IN4(g299), .IN5(
        n1497), .QN(n1488) );
  OA221X1 U2399 ( .IN1(n583), .IN2(DFF_350_n1), .IN3(n577), .IN4(n1636), .IN5(
        n1498), .Q(n1487) );
  NAND4X0 U2400 ( .IN1(n1514), .IN2(n1515), .IN3(n1516), .IN4(n1517), .QN(
        g10721) );
  OA22X1 U2401 ( .IN1(n577), .IN2(n1652), .IN3(n583), .IN4(DFF_242_n1), .Q(
        n1514) );
  AOI222X1 U2402 ( .IN1(n1485), .IN2(g1574), .IN3(n1482), .IN4(g293), .IN5(
        n1483), .IN6(g269), .QN(n1515) );
  AOI221X1 U2403 ( .IN1(n1479), .IN2(g1555), .IN3(n1480), .IN4(g1598), .IN5(
        n1522), .QN(n1516) );
  NAND4X0 U2404 ( .IN1(n1533), .IN2(n1534), .IN3(n1535), .IN4(n1536), .QN(
        g10719) );
  AOI222X1 U2405 ( .IN1(n1479), .IN2(g1549), .IN3(n572), .IN4(g1744), .IN5(
        n1480), .IN6(g1592), .QN(n1533) );
  OA221X1 U2406 ( .IN1(n583), .IN2(DFF_168_n1), .IN3(n577), .IN4(n1649), .IN5(
        n1549), .Q(n1535) );
  NAND4X0 U2407 ( .IN1(n1468), .IN2(n1469), .IN3(n1470), .IN4(n1471), .QN(
        g10726) );
  AOI222X1 U2408 ( .IN1(n1479), .IN2(g1564), .IN3(n572), .IN4(g1759), .IN5(
        n1480), .IN6(g1607), .QN(n1470) );
  AOI222X1 U2409 ( .IN1(n1484), .IN2(n1650), .IN3(n1485), .IN4(g1583), .IN5(
        n1486), .IN6(g1540), .QN(n1468) );
  OA221X1 U2410 ( .IN1(n1472), .IN2(n1638), .IN3(n1491), .IN4(n1492), .IN5(
        n1493), .Q(n1490) );
  NAND2X0 U2411 ( .IN1(n573), .IN2(n1477), .QN(n1492) );
  OA221X1 U2412 ( .IN1(n1472), .IN2(n1639), .IN3(n1473), .IN4(n1474), .IN5(
        n1475), .Q(n1471) );
  NAND2X0 U2413 ( .IN1(n1477), .IN2(n1478), .QN(n1474) );
  AO222X1 U2414 ( .IN1(n572), .IN2(g1750), .IN3(n579), .IN4(g9), .IN5(n575), 
        .IN6(g1727), .Q(n1522) );
  AO222X1 U2415 ( .IN1(g1333), .IN2(n576), .IN3(g1308), .IN4(n1511), .IN5(
        g4214), .IN6(n1476), .Q(n1562) );
  AO22X1 U2416 ( .IN1(n1480), .IN2(g1604), .IN3(n1479), .IN4(g1561), .Q(n1497)
         );
  AO22X1 U2417 ( .IN1(g4202), .IN2(n1481), .IN3(g944), .IN4(n1506), .Q(n1563)
         );
  ISOLANDX1 U2418 ( .D(g968), .ISO(n1472), .Q(n1564) );
  NOR4X0 U2419 ( .IN1(n1537), .IN2(n1538), .IN3(n1539), .IN4(n1540), .QN(n1536) );
  AO222X1 U2420 ( .IN1(g950), .IN2(n580), .IN3(g928), .IN4(n1508), .IN5(g971), 
        .IN6(n1506), .Q(n1539) );
  AO222X1 U2421 ( .IN1(g4204), .IN2(n1530), .IN3(g119), .IN4(n579), .IN5(g4191), .IN6(n1507), .Q(n1538) );
  NAND3X0 U2422 ( .IN1(n574), .IN2(n1541), .IN3(n1542), .QN(n1537) );
  NAND2X0 U2423 ( .IN1(g123), .IN2(n578), .QN(n1542) );
  INVX0 U2424 ( .IN(n1509), .QN(n574) );
  NOR3X0 U2425 ( .IN1(n1518), .IN2(n1519), .IN3(n1520), .QN(n1517) );
  AO222X1 U2426 ( .IN1(g981), .IN2(n1506), .IN3(g956), .IN4(n580), .IN5(g4198), 
        .IN6(n1481), .Q(n1520) );
  AOI22X1 U2427 ( .IN1(g4200), .IN2(n1481), .IN3(g1580), .IN4(n1485), .QN(
        n1498) );
  AOI22X1 U2428 ( .IN1(n575), .IN2(g1733), .IN3(n572), .IN4(g1756), .QN(n1496)
         );
  AOI222X1 U2429 ( .IN1(n1485), .IN2(g1567), .IN3(n1482), .IN4(g287), .IN5(
        n1483), .IN6(g263), .QN(n1549) );
  OA22X1 U2430 ( .IN1(n1543), .IN2(n1568), .IN3(n1550), .IN4(n1640), .Q(n1559)
         );
  NAND2X0 U2431 ( .IN1(n573), .IN2(n1478), .QN(n1568) );
  NAND2X0 U2432 ( .IN1(g1317), .IN2(n550), .QN(n1255) );
  NAND3X0 U2433 ( .IN1(n1113), .IN2(n1270), .IN3(n629), .QN(n1227) );
  NAND4X0 U2434 ( .IN1(n1271), .IN2(n1272), .IN3(n1273), .IN4(n1274), .QN(
        n1270) );
  XNOR2X1 U2435 ( .IN1(test_so2), .IN2(g1255), .Q(n1271) );
  XNOR2X1 U2436 ( .IN1(g1015), .IN2(g1265), .Q(n1272) );
  AO21X1 U2437 ( .IN1(g201), .IN2(n1880), .IN3(n1288), .Q(n1261) );
  OA221X1 U2438 ( .IN1(n1289), .IN2(n1699), .IN3(n627), .IN4(n1290), .IN5(
        n1959), .Q(n1288) );
  INVX0 U2439 ( .IN(n1289), .QN(n627) );
  AO22X1 U2440 ( .IN1(g1766), .IN2(n1653), .IN3(n1882), .IN4(g10719), .Q(n1373) );
  AO22X1 U2441 ( .IN1(g1776), .IN2(n1653), .IN3(n1882), .IN4(g10721), .Q(n1374) );
  AO22X1 U2442 ( .IN1(n1862), .IN2(n1863), .IN3(n1864), .IN4(g1280), .Q(n1326)
         );
  OAI21X1 U2443 ( .IN1(n1328), .IN2(n1329), .IN3(n1864), .QN(n1863) );
  INVX0 U2444 ( .IN(g109), .QN(n1988) );
  INVX0 U2445 ( .IN(g109), .QN(n1987) );
  AO22X1 U2446 ( .IN1(n549), .IN2(g1791), .IN3(g1324), .IN4(n1255), .Q(g11607)
         );
  AO22X1 U2447 ( .IN1(n549), .IN2(g1776), .IN3(g1314), .IN4(n1255), .Q(g11604)
         );
  AO22X1 U2448 ( .IN1(n549), .IN2(g1781), .IN3(g1318), .IN4(n1255), .Q(g11605)
         );
  AO22X1 U2449 ( .IN1(n549), .IN2(g1796), .IN3(g1327), .IN4(n1255), .Q(g11608)
         );
  AO22X1 U2450 ( .IN1(n549), .IN2(g1786), .IN3(g1321), .IN4(n1255), .Q(g11606)
         );
  AO22X1 U2451 ( .IN1(g546), .IN2(n1925), .IN3(n1954), .IN4(n1412), .Q(g10791)
         );
  AO22X1 U2452 ( .IN1(g575), .IN2(n1927), .IN3(n1954), .IN4(n1411), .Q(g10800)
         );
  AO22X1 U2453 ( .IN1(g557), .IN2(n1926), .IN3(n1954), .IN4(n1408), .Q(g10795)
         );
  AO22X1 U2454 ( .IN1(g549), .IN2(n1927), .IN3(n1954), .IN4(n1409), .Q(g10855)
         );
  AO22X1 U2455 ( .IN1(g1678), .IN2(n1929), .IN3(n1955), .IN4(n1408), .Q(g10862) );
  AO22X1 U2456 ( .IN1(g1675), .IN2(n1928), .IN3(n1955), .IN4(n1410), .Q(g10860) );
  AO22X1 U2457 ( .IN1(g554), .IN2(n1926), .IN3(n1954), .IN4(n1410), .Q(g10793)
         );
  AO22X1 U2458 ( .IN1(g1672), .IN2(n1928), .IN3(n1954), .IN4(n1412), .Q(g10858) );
  AO22X1 U2459 ( .IN1(g1666), .IN2(n1888), .IN3(n1406), .IN4(n1875), .Q(g10863) );
  OA21X1 U2460 ( .IN1(n532), .IN2(g1718), .IN3(n1407), .Q(n1406) );
  AO22X1 U2461 ( .IN1(n549), .IN2(test_so5), .IN3(test_so9), .IN4(n1255), .Q(
        g11603) );
  AO22X1 U2462 ( .IN1(n549), .IN2(g1801), .IN3(g1330), .IN4(n1255), .Q(g11609)
         );
  AO22X1 U2463 ( .IN1(n549), .IN2(g1806), .IN3(g1333), .IN4(n1255), .Q(g11610)
         );
  AO22X1 U2464 ( .IN1(n549), .IN2(g1766), .IN3(g1308), .IN4(n1255), .Q(g11602)
         );
  AO22X1 U2465 ( .IN1(g1663), .IN2(n1888), .IN3(n1875), .IN4(n1409), .Q(g10861) );
  AO22X1 U2466 ( .IN1(g1660), .IN2(n1888), .IN3(n1875), .IN4(n1411), .Q(g10859) );
  AO221X1 U2467 ( .IN1(test_so5), .IN2(n1373), .IN3(g1781), .IN4(n1374), .IN5(
        n1881), .Q(n1368) );
  ISOLANDX1 U2468 ( .D(g1336), .ISO(n1227), .Q(n1231) );
  NOR2X0 U2469 ( .IN1(n1223), .IN2(n1224), .QN(g11641) );
  OA22X1 U2470 ( .IN1(n687), .IN2(n1225), .IN3(n1226), .IN4(n1721), .Q(n1223)
         );
  NOR2X0 U2471 ( .IN1(n1227), .IN2(n1228), .QN(n1226) );
  NOR2X0 U2472 ( .IN1(n1233), .IN2(n1224), .QN(g11639) );
  XNOR2X1 U2473 ( .IN1(g1341), .IN2(n1231), .Q(n1233) );
  NOR2X0 U2474 ( .IN1(n1234), .IN2(n1224), .QN(g11636) );
  XOR2X1 U2475 ( .IN1(n1227), .IN2(g1336), .Q(n1234) );
  NOR2X0 U2476 ( .IN1(n1230), .IN2(n1224), .QN(g11640) );
  AOI22X1 U2477 ( .IN1(n1231), .IN2(n1232), .IN3(n1225), .IN4(g1346), .QN(
        n1230) );
  ISOLANDX1 U2478 ( .D(g1341), .ISO(n1229), .Q(n1232) );
  XNOR2X1 U2479 ( .IN1(n1332), .IN2(g1027), .Q(n1285) );
  NAND2X0 U2480 ( .IN1(g1032), .IN2(n1222), .QN(n1332) );
  NOR3X0 U2481 ( .IN1(n1281), .IN2(n1282), .IN3(n1283), .QN(n1273) );
  XOR2X1 U2482 ( .IN1(test_so6), .IN2(g1023), .Q(n1281) );
  XOR2X1 U2483 ( .IN1(g1260), .IN2(g1019), .Q(n1283) );
  XOR2X1 U2484 ( .IN1(n1284), .IN2(n1285), .Q(n1282) );
  AO22X1 U2485 ( .IN1(g1618), .IN2(n1930), .IN3(n1955), .IN4(n1256), .Q(g11579) );
  XOR2X1 U2486 ( .IN1(g1610), .IN2(n1257), .Q(n1256) );
  OA22X1 U2487 ( .IN1(n1258), .IN2(n1259), .IN3(n1260), .IN4(n1261), .Q(n1257)
         );
  ISOLANDX1 U2488 ( .D(n1262), .ISO(n1258), .Q(n1260) );
  OAI22X1 U2489 ( .IN1(n1375), .IN2(n715), .IN3(n1032), .IN4(n1376), .QN(
        g11293) );
  OA21X1 U2490 ( .IN1(n1377), .IN2(DFF_311_n1), .IN3(n815), .Q(n1376) );
  OA22X1 U2491 ( .IN1(g10719), .IN2(n1653), .IN3(g1806), .IN4(n1882), .Q(n1375) );
  AND3X1 U2492 ( .IN1(n1378), .IN2(n1379), .IN3(g4904), .Q(n1377) );
  AND3X1 U2493 ( .IN1(n1956), .IN2(n1610), .IN3(g1289), .Q(n1113) );
  INVX0 U2494 ( .IN(n1924), .QN(n1956) );
  NOR3X0 U2495 ( .IN1(n1983), .IN2(n1865), .IN3(n1866), .QN(n1362) );
  NAND3X0 U2496 ( .IN1(n1977), .IN2(DFF_121_n1), .IN3(g2986), .QN(n1059) );
  NAND3X0 U2497 ( .IN1(n1977), .IN2(DFF_194_n1), .IN3(g3069), .QN(n1236) );
  AO22X1 U2498 ( .IN1(g1796), .IN2(n1653), .IN3(n1882), .IN4(g10663), .Q(n1372) );
  AO22X1 U2499 ( .IN1(g1786), .IN2(n1653), .IN3(n1882), .IN4(g10724), .Q(n1371) );
  OR2X1 U2500 ( .IN1(n1484), .IN2(g6254), .Q(n1867) );
  AO22X1 U2501 ( .IN1(g1275), .IN2(n1113), .IN3(g1235), .IN4(n1120), .Q(g7296)
         );
  AO22X1 U2502 ( .IN1(g1304), .IN2(n1113), .IN3(g1300), .IN4(n1120), .Q(g7291)
         );
  AO22X1 U2503 ( .IN1(g1292), .IN2(n1113), .IN3(g1284), .IN4(n1120), .Q(g7294)
         );
  AO22X1 U2504 ( .IN1(g1255), .IN2(n1113), .IN3(g1260), .IN4(n1120), .Q(g7301)
         );
  AO22X1 U2505 ( .IN1(g1284), .IN2(n1113), .IN3(g1280), .IN4(n1120), .Q(g7295)
         );
  AO22X1 U2506 ( .IN1(g1250), .IN2(n1113), .IN3(g1255), .IN4(n1120), .Q(g7300)
         );
  AO22X1 U2507 ( .IN1(g1240), .IN2(n1113), .IN3(g1245), .IN4(n1120), .Q(g7298)
         );
  AO22X1 U2508 ( .IN1(g1265), .IN2(n1113), .IN3(test_so6), .IN4(n1120), .Q(
        g7303) );
  AO22X1 U2509 ( .IN1(g1296), .IN2(n1113), .IN3(g1292), .IN4(n1120), .Q(g7293)
         );
  AO22X1 U2510 ( .IN1(g1245), .IN2(n1113), .IN3(g1250), .IN4(n1120), .Q(g7299)
         );
  AO22X1 U2511 ( .IN1(g1235), .IN2(n1113), .IN3(g1240), .IN4(n1120), .Q(g7297)
         );
  AO22X1 U2512 ( .IN1(g1300), .IN2(n1113), .IN3(g1296), .IN4(n1120), .Q(g7292)
         );
  AO22X1 U2513 ( .IN1(g1260), .IN2(n1113), .IN3(g1265), .IN4(n1120), .Q(g7302)
         );
  AO22X1 U2514 ( .IN1(test_so6), .IN2(n1113), .IN3(g1304), .IN4(n1120), .Q(
        g7290) );
  AO22X1 U2515 ( .IN1(g105), .IN2(n1930), .IN3(n1955), .IN4(n1393), .Q(g10898)
         );
  NAND2X0 U2516 ( .IN1(n1394), .IN2(n1222), .QN(n1393) );
  XOR3X1 U2517 ( .IN1(n1397), .IN2(n1398), .IN3(n1399), .Q(n1394) );
  XNOR2X1 U2518 ( .IN1(g1023), .IN2(g1027), .Q(n1399) );
  AO22X1 U2519 ( .IN1(n1875), .IN2(n1453), .IN3(g1654), .IN4(n1888), .Q(g10765) );
  AO22X1 U2520 ( .IN1(g1724), .IN2(n1451), .IN3(n528), .IN4(n561), .Q(g10771)
         );
  INVX0 U2521 ( .IN(n1414), .QN(n528) );
  AO22X1 U2522 ( .IN1(n1113), .IN2(n1284), .IN3(g1275), .IN4(n1120), .Q(g11443) );
  AO22X1 U2523 ( .IN1(g569), .IN2(n1928), .IN3(n1955), .IN4(n1453), .Q(g10717)
         );
  AO22X1 U2524 ( .IN1(g1687), .IN2(n1925), .IN3(n1954), .IN4(n1417), .Q(g10776) );
  AO22X1 U2525 ( .IN1(g566), .IN2(n1927), .IN3(n1954), .IN4(n1417), .Q(g10799)
         );
  AO22X1 U2526 ( .IN1(g563), .IN2(n1927), .IN3(n1954), .IN4(n1402), .Q(g10798)
         );
  AO22X1 U2527 ( .IN1(g1684), .IN2(n1929), .IN3(n1955), .IN4(n1402), .Q(g10866) );
  AO22X1 U2528 ( .IN1(g1733), .IN2(n1451), .IN3(n561), .IN4(n1382), .Q(g10711)
         );
  AO22X1 U2529 ( .IN1(n561), .IN2(n532), .IN3(g1727), .IN4(n1451), .Q(g10773)
         );
  AO22X1 U2530 ( .IN1(n561), .IN2(n534), .IN3(g1721), .IN4(n1451), .Q(g10770)
         );
  AO221X1 U2531 ( .IN1(g1791), .IN2(n1371), .IN3(g1801), .IN4(n1372), .IN5(
        n1882), .Q(n1370) );
  NOR2X0 U2532 ( .IN1(n1868), .IN2(n1967), .QN(n1363) );
  ISOLANDX1 U2533 ( .D(g178), .ISO(n1966), .Q(g6786) );
  ISOLANDX1 U2534 ( .D(g1424), .ISO(n1967), .Q(g6234) );
  AO21X1 U2535 ( .IN1(g123), .IN2(n1968), .IN3(n1132), .Q(g7032) );
  NOR4X0 U2536 ( .IN1(n1133), .IN2(n1134), .IN3(n1135), .IN4(n1136), .QN(n1132) );
  OR4X1 U2537 ( .IN1(g148), .IN2(g153), .IN3(g158), .IN4(g162), .Q(n1133) );
  OR4X1 U2538 ( .IN1(g131), .IN2(g135), .IN3(g139), .IN4(g143), .Q(n1134) );
  INVX0 U2539 ( .IN(g1703), .QN(n744) );
  OA21X1 U2540 ( .IN1(n1107), .IN2(n1108), .IN3(n1109), .Q(g7586) );
  OA21X1 U2541 ( .IN1(n1110), .IN2(n1103), .IN3(g1227), .Q(n1108) );
  AND4X1 U2542 ( .IN1(n1110), .IN2(g1218), .IN3(g1223), .IN4(n557), .Q(n1107)
         );
  NOR2X0 U2543 ( .IN1(n1965), .IN2(n1286), .QN(g11514) );
  XOR3X1 U2544 ( .IN1(n1261), .IN2(g1415), .IN3(n1287), .Q(n1286) );
  XOR3X1 U2545 ( .IN1(g1515), .IN2(g1448), .IN3(n1602), .Q(n1287) );
  AO22X1 U2546 ( .IN1(g1), .IN2(n1975), .IN3(n1154), .IN4(n1155), .Q(g6679) );
  NOR2X0 U2547 ( .IN1(n1156), .IN2(n1157), .QN(n1155) );
  NOR4X0 U2548 ( .IN1(n1158), .IN2(n1710), .IN3(n1602), .IN4(n1627), .QN(n1154) );
  OR4X1 U2549 ( .IN1(g1403), .IN2(g1407), .IN3(g1411), .IN4(g1415), .Q(n1156)
         );
  XNOR2X1 U2550 ( .IN1(n1381), .IN2(n1382), .Q(n1378) );
  OA22X1 U2551 ( .IN1(g1857), .IN2(n1380), .IN3(n1682), .IN4(n920), .Q(n1381)
         );
  OR2X1 U2552 ( .IN1(g845), .IN2(g849), .Q(n1443) );
  NAND4X0 U2553 ( .IN1(g6234), .IN2(n1159), .IN3(g1432), .IN4(g1448), .QN(
        n1158) );
  NOR2X0 U2554 ( .IN1(n1111), .IN2(n540), .QN(g7581) );
  XOR2X1 U2555 ( .IN1(n1112), .IN2(g1223), .Q(n1111) );
  NAND2X0 U2556 ( .IN1(n557), .IN2(g1218), .QN(n1112) );
  NOR2X0 U2557 ( .IN1(n1102), .IN2(n540), .QN(g7632) );
  XOR2X1 U2558 ( .IN1(n1103), .IN2(g1218), .Q(n1102) );
  NAND4X0 U2559 ( .IN1(g182), .IN2(g6786), .IN3(n1137), .IN4(g166), .QN(n1136)
         );
  NOR2X0 U2560 ( .IN1(n1106), .IN2(n540), .QN(g7590) );
  AOI21X1 U2561 ( .IN1(n665), .IN2(n557), .IN3(g1231), .QN(n1106) );
  INVX0 U2562 ( .IN(n1724), .QN(n560) );
  AO22X1 U2563 ( .IN1(g1687), .IN2(n1882), .IN3(g1669), .IN4(n1653), .Q(g6955)
         );
  AO22X1 U2564 ( .IN1(g1684), .IN2(n1882), .IN3(g1666), .IN4(n1653), .Q(g6949)
         );
  AO22X1 U2565 ( .IN1(g1681), .IN2(n1882), .IN3(g1663), .IN4(n1653), .Q(g6942)
         );
  AO22X1 U2566 ( .IN1(g1678), .IN2(n1882), .IN3(g1660), .IN4(n1653), .Q(g6932)
         );
  AO22X1 U2567 ( .IN1(g1675), .IN2(n1882), .IN3(g1657), .IN4(n1653), .Q(g6926)
         );
  AO22X1 U2568 ( .IN1(g1672), .IN2(n1882), .IN3(g1654), .IN4(n1653), .Q(g6920)
         );
  AO21X1 U2569 ( .IN1(g617), .IN2(n959), .IN3(n960), .Q(n899) );
  AO21X1 U2570 ( .IN1(g1840), .IN2(n926), .IN3(n929), .Q(n853) );
  NAND4X0 U2571 ( .IN1(n1184), .IN2(n1185), .IN3(n1186), .IN4(n1187), .QN(
        n1183) );
  NOR4X0 U2572 ( .IN1(n1188), .IN2(g192), .IN3(g248), .IN4(g197), .QN(n1187)
         );
  AND3X1 U2573 ( .IN1(n1977), .IN2(n1700), .IN3(g201), .Q(n1186) );
  NAND3X0 U2574 ( .IN1(n1711), .IN2(n1629), .IN3(n1603), .QN(n1188) );
  NAND2X0 U2575 ( .IN1(g1765), .IN2(g1610), .QN(n1217) );
  NAND2X0 U2576 ( .IN1(n1137), .IN2(n1613), .QN(n1145) );
  NOR2X0 U2577 ( .IN1(n1964), .IN2(test_so1), .QN(n1046) );
  NOR2X0 U2578 ( .IN1(n1724), .IN2(g4089), .QN(g6842) );
  AO22X1 U2579 ( .IN1(g673), .IN2(n899), .IN3(n648), .IN4(n914), .Q(n913) );
  XOR2X1 U2580 ( .IN1(g658), .IN2(n718), .Q(n914) );
  AO22X1 U2581 ( .IN1(g1887), .IN2(n853), .IN3(n622), .IN4(n871), .Q(n870) );
  XOR2X1 U2582 ( .IN1(g1872), .IN2(n712), .Q(n871) );
  NOR2X0 U2583 ( .IN1(n892), .IN2(g1891), .QN(n877) );
  NOR2X0 U2584 ( .IN1(n950), .IN2(g677), .QN(n935) );
  NAND2X0 U2585 ( .IN1(g1104), .IN2(n985), .QN(n978) );
  NAND2X0 U2586 ( .IN1(g461), .IN2(n1641), .QN(n1306) );
  NOR2X0 U2587 ( .IN1(n662), .IN2(g1718), .QN(n1404) );
  OA21X1 U2588 ( .IN1(n1609), .IN2(g591), .IN3(n668), .Q(n1160) );
  OA21X1 U2589 ( .IN1(n1655), .IN2(g1814), .IN3(n715), .Q(n1148) );
  NAND2X0 U2590 ( .IN1(g599), .IN2(n1593), .QN(n953) );
  NAND2X0 U2591 ( .IN1(g599), .IN2(n1607), .QN(n1025) );
  NAND2X0 U2592 ( .IN1(g1822), .IN2(n1608), .QN(n920) );
  AO21X1 U2593 ( .IN1(g869), .IN2(n1352), .IN3(n1966), .Q(n1334) );
  NAND2X0 U2594 ( .IN1(n1724), .IN2(n744), .QN(n1054) );
  NAND2X0 U2595 ( .IN1(n1970), .IN2(DFF_441_n1), .QN(n1345) );
  NOR2X0 U2596 ( .IN1(n1965), .IN2(g869), .QN(n1384) );
  AND3X1 U2597 ( .IN1(g743), .IN2(n1969), .IN3(g744), .Q(g5659) );
  AND3X1 U2598 ( .IN1(g741), .IN2(n1976), .IN3(g742), .Q(g5658) );
  NAND2X0 U2599 ( .IN1(g4180), .IN2(n1093), .QN(n1092) );
  NAND2X0 U2600 ( .IN1(g466), .IN2(n1606), .QN(n1307) );
  NOR3X0 U2601 ( .IN1(g591), .IN2(g611), .IN3(n964), .QN(n954) );
  NAND2X0 U2602 ( .IN1(g471), .IN2(n1646), .QN(n1325) );
  NOR2X0 U2603 ( .IN1(n1962), .IN2(g1212), .QN(n1109) );
  NAND2X0 U2604 ( .IN1(g591), .IN2(n1644), .QN(n966) );
  NAND2X0 U2605 ( .IN1(g627), .IN2(n1612), .QN(n1119) );
  NOR2X0 U2606 ( .IN1(n1966), .IN2(g1718), .QN(n1416) );
  NOR4X0 U2607 ( .IN1(n1654), .IN2(g1104), .IN3(g1107), .IN4(g1110), .QN(n1263) );
  NOR2X0 U2608 ( .IN1(n1614), .IN2(g1110), .QN(n985) );
  NAND3X0 U2609 ( .IN1(g745), .IN2(n1976), .IN3(g746), .QN(n1042) );
  NOR3X0 U2610 ( .IN1(g1814), .IN2(g1834), .IN3(n928), .QN(n1032) );
  NAND2X0 U2611 ( .IN1(g1231), .IN2(n665), .QN(n1114) );
  NAND3X0 U2612 ( .IN1(n1884), .IN2(g461), .IN3(g466), .QN(n1302) );
  NAND3X0 U2613 ( .IN1(n1614), .IN2(n1677), .IN3(g1104), .QN(n993) );
  NAND3X0 U2614 ( .IN1(n1646), .IN2(n1606), .IN3(g461), .QN(n1318) );
  NAND3X0 U2615 ( .IN1(test_so5), .IN2(g1766), .IN3(g1776), .QN(n1172) );
  NAND3X0 U2616 ( .IN1(n1658), .IN2(n1614), .IN3(g1110), .QN(n999) );
  NAND2X0 U2617 ( .IN1(g219), .IN2(g2355), .QN(n974) );
  NAND2X0 U2618 ( .IN1(g231), .IN2(g2355), .QN(n995) );
  NAND2X0 U2619 ( .IN1(g207), .IN2(g2355), .QN(n1001) );
  NAND2X0 U2620 ( .IN1(g225), .IN2(n1880), .QN(n981) );
  NAND2X0 U2621 ( .IN1(g186), .IN2(n1880), .QN(n989) );
  NAND2X0 U2622 ( .IN1(g237), .IN2(n1880), .QN(n1007) );
  NAND2X0 U2623 ( .IN1(g213), .IN2(n1880), .QN(n1012) );
  NAND2X0 U2624 ( .IN1(g1504), .IN2(n1969), .QN(n1166) );
  NAND2X0 U2625 ( .IN1(n1969), .IN2(DFF_126_n1), .QN(n1216) );
  NAND2X0 U2626 ( .IN1(g4174), .IN2(g4173), .QN(n1214) );
  NOR3X0 U2627 ( .IN1(g650), .IN2(g654), .IN3(n1128), .QN(n959) );
  NAND2X0 U2628 ( .IN1(g1828), .IN2(g1814), .QN(n817) );
  AND4X1 U2629 ( .IN1(n1845), .IN2(n1843), .IN3(n1847), .IN4(n799), .Q(n795)
         );
  NOR2X0 U2630 ( .IN1(g6258), .IN2(g6257), .QN(n799) );
  AO21X1 U2631 ( .IN1(n605), .IN2(n930), .IN3(n606), .Q(g8920) );
  XNOR2X1 U2632 ( .IN1(g713), .IN2(n931), .Q(n930) );
  NAND2X0 U2633 ( .IN1(n850), .IN2(n932), .QN(n931) );
  AO222X1 U2634 ( .IN1(n933), .IN2(n934), .IN3(n935), .IN4(n936), .IN5(g718), 
        .IN6(n899), .Q(n932) );
  NAND2X0 U2635 ( .IN1(g1814), .IN2(n1643), .QN(n826) );
  NAND2X0 U2636 ( .IN1(g1822), .IN2(n1605), .QN(n822) );
  NAND2X0 U2637 ( .IN1(g668), .IN2(n913), .QN(n912) );
  NAND2X0 U2638 ( .IN1(g1882), .IN2(n870), .QN(n869) );
  ISOLANDX1 U2639 ( .D(n962), .ISO(n958), .Q(n804) );
  OAI22X1 U2640 ( .IN1(n1696), .IN2(n902), .IN3(n901), .IN4(g731), .QN(n962)
         );
  ISOLANDX1 U2641 ( .D(n1147), .ISO(g1868), .Q(n926) );
  NAND3X0 U2642 ( .IN1(g1223), .IN2(g1218), .IN3(g1227), .QN(n1110) );
  NAND3X0 U2643 ( .IN1(n1607), .IN2(n1644), .IN3(g605), .QN(n832) );
  AND4X1 U2644 ( .IN1(n1624), .IN2(n1687), .IN3(n1206), .IN4(n1207), .Q(n1185)
         );
  NOR2X0 U2645 ( .IN1(g1386), .IN2(g1383), .QN(n1206) );
  NOR4X0 U2646 ( .IN1(g219), .IN2(g213), .IN3(g207), .IN4(g186), .QN(n1207) );
  NAND2X0 U2647 ( .IN1(g4176), .IN2(n1193), .QN(n1153) );
  NAND2X0 U2648 ( .IN1(g4178), .IN2(n1125), .QN(n1099) );
  AND4X1 U2649 ( .IN1(n936), .IN2(n1615), .IN3(n965), .IN4(n1662), .Q(n907) );
  NOR2X0 U2650 ( .IN1(g713), .IN2(g677), .QN(n965) );
  AND4X1 U2651 ( .IN1(n878), .IN2(n1616), .IN3(n919), .IN4(n1663), .Q(n862) );
  NOR2X0 U2652 ( .IN1(g1927), .IN2(g1891), .QN(n919) );
  NAND2X0 U2653 ( .IN1(g798), .IN2(g794), .QN(n1029) );
  ISOLANDX1 U2654 ( .D(g746), .ISO(g750), .Q(g4171) );
  NAND3X0 U2655 ( .IN1(n959), .IN2(n1609), .IN3(g617), .QN(n1016) );
  NAND3X0 U2656 ( .IN1(n926), .IN2(n1655), .IN3(g1840), .QN(n1031) );
  NOR2X0 U2657 ( .IN1(g611), .IN2(n834), .QN(n1024) );
  ISOLANDX1 U2658 ( .D(n917), .ISO(n918), .Q(n812) );
  OAI22X1 U2659 ( .IN1(n1697), .IN2(n857), .IN3(n856), .IN4(g1945), .QN(n917)
         );
  AND3X1 U2660 ( .IN1(g1909), .IN2(g1900), .IN3(g1918), .Q(n876) );
  AND3X1 U2661 ( .IN1(g695), .IN2(g686), .IN3(g704), .Q(n934) );
  NAND2X0 U2662 ( .IN1(n1007), .IN2(n1008), .QN(n969) );
  AO221X1 U2663 ( .IN1(n1009), .IN2(g1145), .IN3(n1617), .IN4(n1010), .IN5(
        g2355), .Q(n1008) );
  NOR2X0 U2664 ( .IN1(n999), .IN2(n1654), .QN(n1009) );
  NAND2X0 U2665 ( .IN1(g1101), .IN2(n634), .QN(n1010) );
  NAND2X0 U2666 ( .IN1(n1012), .IN2(n1013), .QN(n979) );
  AO221X1 U2667 ( .IN1(n1014), .IN2(g1129), .IN3(n1705), .IN4(n1015), .IN5(
        n1880), .Q(n1013) );
  NAND2X0 U2668 ( .IN1(n633), .IN2(g1101), .QN(n1015) );
  NOR2X0 U2669 ( .IN1(n1654), .IN2(n1005), .QN(n1014) );
  NAND2X0 U2670 ( .IN1(n1001), .IN2(n1002), .QN(n986) );
  AO221X1 U2671 ( .IN1(n1003), .IN2(g1125), .IN3(n1708), .IN4(n1004), .IN5(
        n1880), .Q(n1002) );
  NAND2X0 U2672 ( .IN1(n633), .IN2(n1654), .QN(n1004) );
  NOR2X0 U2673 ( .IN1(g1101), .IN2(n1005), .QN(n1003) );
  NAND2X0 U2674 ( .IN1(n974), .IN2(n975), .QN(n973) );
  AO221X1 U2675 ( .IN1(n976), .IN2(g1133), .IN3(n1706), .IN4(n977), .IN5(n1880), .Q(n975) );
  NAND2X0 U2676 ( .IN1(n631), .IN2(n1654), .QN(n977) );
  NOR2X0 U2677 ( .IN1(g1101), .IN2(n978), .QN(n976) );
  NOR2X0 U2678 ( .IN1(g4173), .IN2(n537), .QN(g4940) );
  NAND2X0 U2679 ( .IN1(g4181), .IN2(n630), .QN(n1045) );
  AO22X1 U2680 ( .IN1(g192), .IN2(n1880), .IN3(g1512), .IN4(n1959), .Q(n1082)
         );
  AO22X1 U2681 ( .IN1(g243), .IN2(n1880), .IN3(g1633), .IN4(n1959), .Q(n1069)
         );
  AO22X1 U2682 ( .IN1(g248), .IN2(g2355), .IN3(g1636), .IN4(n1959), .Q(n1077)
         );
  ISOLANDX1 U2683 ( .D(g382), .ISO(n1385), .Q(n1420) );
  AO22X1 U2684 ( .IN1(g192), .IN2(g2355), .IN3(g549), .IN4(n1959), .Q(g6049)
         );
  AO22X1 U2685 ( .IN1(g248), .IN2(n1880), .IN3(g575), .IN4(n1959), .Q(g6045)
         );
  AO22X1 U2686 ( .IN1(g243), .IN2(g2355), .IN3(g572), .IN4(n1959), .Q(g6042)
         );
  AO21X1 U2687 ( .IN1(n805), .IN2(n963), .IN3(n649), .Q(n958) );
  NAND2X0 U2688 ( .IN1(g639), .IN2(n964), .QN(n963) );
  NAND4X0 U2689 ( .IN1(n648), .IN2(g668), .IN3(g658), .IN4(n908), .QN(n949) );
  NAND4X0 U2690 ( .IN1(n622), .IN2(g1882), .IN3(g1872), .IN4(n863), .QN(n891)
         );
  AO21X1 U2691 ( .IN1(g1639), .IN2(n1922), .IN3(n1049), .Q(g8193) );
  OA221X1 U2692 ( .IN1(n1050), .IN2(test_so4), .IN3(n1661), .IN4(n1051), .IN5(
        n1953), .Q(n1049) );
  NAND2X0 U2693 ( .IN1(n632), .IN2(n1654), .QN(n1051) );
  NOR2X0 U2694 ( .IN1(g1101), .IN2(n993), .QN(n1050) );
  AND3X1 U2695 ( .IN1(n831), .IN2(n832), .IN3(n833), .Q(n829) );
  NAND2X0 U2696 ( .IN1(n834), .IN2(g599), .QN(n833) );
  OA221X1 U2697 ( .IN1(n806), .IN2(g1834), .IN3(n623), .IN4(n807), .IN5(g2355), 
        .Q(g9555) );
  NAND2X0 U2698 ( .IN1(g1834), .IN2(n808), .QN(n807) );
  ISOLANDX1 U2699 ( .D(n808), .ISO(n623), .Q(n806) );
  AO21X1 U2700 ( .IN1(n809), .IN2(n598), .IN3(g1840), .Q(n808) );
  AND3X1 U2701 ( .IN1(n1044), .IN2(n1045), .IN3(n1046), .Q(g8244) );
  OR2X1 U2702 ( .IN1(g4181), .IN2(n630), .Q(n1044) );
  AND3X1 U2703 ( .IN1(n1215), .IN2(n1214), .IN3(n1046), .Q(g5529) );
  OR2X1 U2704 ( .IN1(g4173), .IN2(g4174), .Q(n1215) );
  AND3X1 U2705 ( .IN1(n1192), .IN2(n1153), .IN3(n1046), .Q(g6123) );
  OR2X1 U2706 ( .IN1(g4176), .IN2(n1193), .Q(n1192) );
  AND3X1 U2707 ( .IN1(n1124), .IN2(n1099), .IN3(n1046), .Q(g7191) );
  OR2X1 U2708 ( .IN1(g4178), .IN2(n1125), .Q(n1124) );
  AND3X1 U2709 ( .IN1(n1091), .IN2(n1092), .IN3(n1046), .Q(g8019) );
  OR2X1 U2710 ( .IN1(n1093), .IN2(g4180), .Q(n1091) );
  AND3X1 U2711 ( .IN1(n1122), .IN2(n1097), .IN3(n520), .Q(g7202) );
  OR2X1 U2712 ( .IN1(g814), .IN2(n1123), .Q(n1122) );
  AND3X1 U2713 ( .IN1(n1190), .IN2(n1151), .IN3(n520), .Q(g6126) );
  OR2X1 U2714 ( .IN1(g806), .IN2(n1191), .Q(n1190) );
  AND3X1 U2715 ( .IN1(n1089), .IN2(n1043), .IN3(n520), .Q(g8024) );
  OR2X1 U2716 ( .IN1(n1090), .IN2(g822), .Q(n1089) );
  AND3X1 U2717 ( .IN1(n1149), .IN2(n1634), .IN3(n1977), .Q(g6747) );
  NAND2X0 U2718 ( .IN1(n1714), .IN2(DFF_452_n1), .QN(n1149) );
  NOR4X0 U2719 ( .IN1(n1203), .IN2(n1204), .IN3(g192), .IN4(g1400), .QN(n1202)
         );
  NAND3X0 U2720 ( .IN1(n1619), .IN2(n1598), .IN3(n1678), .QN(n1204) );
  NAND4X0 U2721 ( .IN1(n1184), .IN2(n1185), .IN3(n1205), .IN4(n1700), .QN(
        n1203) );
  NOR2X0 U2722 ( .IN1(g1397), .IN2(g1389), .QN(n1205) );
  NAND3X0 U2723 ( .IN1(g1786), .IN2(n1141), .IN3(g1791), .QN(n1117) );
  OAI22X1 U2724 ( .IN1(g1153), .IN2(n1685), .IN3(g1149), .IN4(n1265), .QN(
        n1264) );
  OA21X1 U2725 ( .IN1(n1266), .IN2(n1267), .IN3(n1686), .Q(n1265) );
  NAND4X0 U2726 ( .IN1(n1660), .IN2(n1617), .IN3(n1597), .IN4(n1269), .QN(
        n1266) );
  NAND4X0 U2727 ( .IN1(n1661), .IN2(n1618), .IN3(n1596), .IN4(n1268), .QN(
        n1267) );
  OR4X1 U2728 ( .IN1(n826), .IN2(g1828), .IN3(g1834), .IN4(g1840), .Q(n1038)
         );
  NAND2X0 U2729 ( .IN1(n926), .IN2(n927), .QN(n918) );
  AO21X1 U2730 ( .IN1(g1857), .IN2(n928), .IN3(n809), .Q(n927) );
  NAND3X0 U2731 ( .IN1(n1608), .IN2(n1643), .IN3(g1828), .QN(n815) );
  AO21X1 U2732 ( .IN1(g1627), .IN2(n1959), .IN3(n568), .Q(n1086) );
  AO21X1 U2733 ( .IN1(g1630), .IN2(n1958), .IN3(n569), .Q(n1088) );
  AO22X1 U2734 ( .IN1(g1415), .IN2(n1169), .IN3(n538), .IN4(g1567), .Q(g6468)
         );
  AO22X1 U2735 ( .IN1(g1466), .IN2(n1167), .IN3(n539), .IN4(g1555), .Q(g6534)
         );
  AO22X1 U2736 ( .IN1(g1504), .IN2(n1167), .IN3(n539), .IN4(g1528), .Q(g6522)
         );
  AO22X1 U2737 ( .IN1(g1448), .IN2(n1169), .IN3(n538), .IN4(g1607), .Q(g6515)
         );
  AO22X1 U2738 ( .IN1(g1407), .IN2(n1169), .IN3(n538), .IN4(g1586), .Q(g6514)
         );
  AO22X1 U2739 ( .IN1(g1470), .IN2(n1167), .IN3(n539), .IN4(g1552), .Q(g6529)
         );
  AO22X1 U2740 ( .IN1(g1436), .IN2(n1169), .IN3(n538), .IN4(g1598), .Q(g6481)
         );
  AO22X1 U2741 ( .IN1(g1474), .IN2(n1167), .IN3(n539), .IN4(g1549), .Q(g6523)
         );
  AO22X1 U2742 ( .IN1(g1490), .IN2(n1167), .IN3(n539), .IN4(g1537), .Q(g6537)
         );
  AO22X1 U2743 ( .IN1(g1432), .IN2(n1169), .IN3(n538), .IN4(g1595), .Q(g6479)
         );
  AO22X1 U2744 ( .IN1(g1419), .IN2(n1169), .IN3(n538), .IN4(g1577), .Q(g6480)
         );
  AO22X1 U2745 ( .IN1(g1508), .IN2(n1167), .IN3(n539), .IN4(g1524), .Q(g6513)
         );
  AO22X1 U2746 ( .IN1(g1403), .IN2(n1169), .IN3(n538), .IN4(g1592), .Q(g6470)
         );
  AO22X1 U2747 ( .IN1(g1486), .IN2(n1167), .IN3(n539), .IN4(g1540), .Q(g6541)
         );
  AO22X1 U2748 ( .IN1(g1478), .IN2(n1167), .IN3(n539), .IN4(g1546), .Q(g6551)
         );
  AO22X1 U2749 ( .IN1(g1458), .IN2(n1167), .IN3(n539), .IN4(g1561), .Q(g6542)
         );
  AO22X1 U2750 ( .IN1(g1424), .IN2(n1169), .IN3(n538), .IN4(g1583), .Q(g6506)
         );
  AO22X1 U2751 ( .IN1(g1440), .IN2(n1169), .IN3(n538), .IN4(g1601), .Q(g6501)
         );
  AO22X1 U2752 ( .IN1(g1499), .IN2(n1167), .IN3(n539), .IN4(g1531), .Q(g6528)
         );
  AO22X1 U2753 ( .IN1(g1520), .IN2(n1169), .IN3(n538), .IN4(g1571), .Q(g6469)
         );
  AO22X1 U2754 ( .IN1(g1428), .IN2(n1169), .IN3(n538), .IN4(g1589), .Q(g6524)
         );
  AO22X1 U2755 ( .IN1(g1453), .IN2(n1167), .IN3(n539), .IN4(g1564), .Q(g6546)
         );
  AO22X1 U2756 ( .IN1(g1444), .IN2(n1169), .IN3(n538), .IN4(g1604), .Q(g6507)
         );
  AO22X1 U2757 ( .IN1(g1494), .IN2(n1167), .IN3(n539), .IN4(g1534), .Q(g6533)
         );
  AO22X1 U2758 ( .IN1(g1482), .IN2(n1167), .IN3(n539), .IN4(g1543), .Q(g6545)
         );
  AO22X1 U2759 ( .IN1(g1411), .IN2(n1169), .IN3(n538), .IN4(g1580), .Q(g6500)
         );
  AO22X1 U2760 ( .IN1(g1515), .IN2(n1169), .IN3(n538), .IN4(g1574), .Q(g6478)
         );
  AO22X1 U2761 ( .IN1(g1462), .IN2(n1167), .IN3(n539), .IN4(g1558), .Q(g6538)
         );
  AO22X1 U2762 ( .IN1(n624), .IN2(g1923), .IN3(n1039), .IN4(g1932), .Q(g8286)
         );
  AO22X1 U2763 ( .IN1(n650), .IN2(g709), .IN3(n1035), .IN4(g718), .Q(g8433) );
  AO22X1 U2764 ( .IN1(g166), .IN2(n1142), .IN3(n517), .IN4(g299), .Q(g6923) );
  AO22X1 U2765 ( .IN1(g178), .IN2(n1142), .IN3(n517), .IN4(g266), .Q(g6900) );
  AO22X1 U2766 ( .IN1(g158), .IN2(n1142), .IN3(n517), .IN4(g275), .Q(g6915) );
  AO22X1 U2767 ( .IN1(g182), .IN2(n1142), .IN3(n517), .IN4(g263), .Q(g6897) );
  AO22X1 U2768 ( .IN1(g153), .IN2(n1142), .IN3(n517), .IN4(g272), .Q(g6910) );
  AO22X1 U2769 ( .IN1(g139), .IN2(n1142), .IN3(n517), .IN4(g296), .Q(g6916) );
  AO22X1 U2770 ( .IN1(g127), .IN2(n1142), .IN3(n517), .IN4(g287), .Q(g6901) );
  AO22X1 U2771 ( .IN1(g131), .IN2(n1142), .IN3(n517), .IN4(g290), .Q(g6907) );
  AO22X1 U2772 ( .IN1(g143), .IN2(n1142), .IN3(n517), .IN4(g302), .Q(g6929) );
  AO22X1 U2773 ( .IN1(g135), .IN2(n1142), .IN3(n517), .IN4(g293), .Q(g6911) );
  AO22X1 U2774 ( .IN1(g148), .IN2(n1142), .IN3(n517), .IN4(g269), .Q(g6906) );
  AO22X1 U2775 ( .IN1(g174), .IN2(n1142), .IN3(n517), .IN4(g281), .Q(g6928) );
  AO22X1 U2776 ( .IN1(g170), .IN2(n1142), .IN3(n517), .IN4(g284), .Q(g6934) );
  AO22X1 U2777 ( .IN1(g162), .IN2(n1142), .IN3(n517), .IN4(g278), .Q(g6922) );
  AO22X1 U2778 ( .IN1(n954), .IN2(n1017), .IN3(n1018), .IN4(n668), .Q(g8631)
         );
  AO221X1 U2779 ( .IN1(n1027), .IN2(n1028), .IN3(n1029), .IN4(n1030), .IN5(
        n1716), .Q(n1017) );
  AO22X1 U2780 ( .IN1(n720), .IN2(n1713), .IN3(g636), .IN4(n1019), .Q(n1018)
         );
  AO22X1 U2781 ( .IN1(n624), .IN2(g1887), .IN3(n1039), .IN4(g1896), .Q(g8282)
         );
  AO22X1 U2782 ( .IN1(n650), .IN2(g673), .IN3(n1035), .IN4(g682), .Q(g8429) );
  AO22X1 U2783 ( .IN1(n650), .IN2(g718), .IN3(g727), .IN4(n1035), .Q(g8434) );
  AO22X1 U2784 ( .IN1(n624), .IN2(g1914), .IN3(n1039), .IN4(g1923), .Q(g8285)
         );
  AO22X1 U2785 ( .IN1(n624), .IN2(g1932), .IN3(g1941), .IN4(n1039), .Q(g8287)
         );
  AO22X1 U2786 ( .IN1(n650), .IN2(g700), .IN3(n1035), .IN4(g709), .Q(g8432) );
  AO22X1 U2787 ( .IN1(g351), .IN2(n1875), .IN3(g1083), .IN4(n1888), .Q(g6068)
         );
  AO22X1 U2788 ( .IN1(g336), .IN2(n1875), .IN3(test_so7), .IN4(n1888), .Q(
        g6054) );
  AO22X1 U2789 ( .IN1(g339), .IN2(n1875), .IN3(g1071), .IN4(n1888), .Q(g5910)
         );
  AO22X1 U2790 ( .IN1(g357), .IN2(n1875), .IN3(g1089), .IN4(n1888), .Q(g6080)
         );
  AO22X1 U2791 ( .IN1(g348), .IN2(n1875), .IN3(g1080), .IN4(n1888), .Q(g6059)
         );
  AO22X1 U2792 ( .IN1(g342), .IN2(n1875), .IN3(g1074), .IN4(n1888), .Q(g6099)
         );
  AO22X1 U2793 ( .IN1(g354), .IN2(n1875), .IN3(g1086), .IN4(n1888), .Q(g6071)
         );
  AO22X1 U2794 ( .IN1(g366), .IN2(n1875), .IN3(g1098), .IN4(n1888), .Q(g6096)
         );
  AO22X1 U2795 ( .IN1(g363), .IN2(n1875), .IN3(g1095), .IN4(n1888), .Q(g6093)
         );
  AO22X1 U2796 ( .IN1(g345), .IN2(n1875), .IN3(g1077), .IN4(n1888), .Q(g5914)
         );
  AO22X1 U2797 ( .IN1(g360), .IN2(n1875), .IN3(g1092), .IN4(n1888), .Q(g6088)
         );
  AO22X1 U2798 ( .IN1(g1621), .IN2(n1931), .IN3(n1955), .IN4(n986), .Q(g8771)
         );
  AO22X1 U2799 ( .IN1(g1630), .IN2(n1933), .IN3(n1955), .IN4(n971), .Q(g8776)
         );
  AO22X1 U2800 ( .IN1(g1615), .IN2(n1931), .IN3(n1955), .IN4(n987), .Q(g8770)
         );
  AO22X1 U2801 ( .IN1(g1512), .IN2(n1931), .IN3(n1955), .IN4(n1047), .Q(g8194)
         );
  XOR2X1 U2802 ( .IN1(n1596), .IN2(n1048), .Q(n1047) );
  NAND4X0 U2803 ( .IN1(g1104), .IN2(g1110), .IN3(n1654), .IN4(n1614), .QN(
        n1048) );
  AO22X1 U2804 ( .IN1(g1636), .IN2(n1924), .IN3(n1954), .IN4(n969), .Q(g8779)
         );
  AO22X1 U2805 ( .IN1(g1624), .IN2(n1932), .IN3(n1955), .IN4(n979), .Q(g8773)
         );
  AO22X1 U2806 ( .IN1(g1627), .IN2(n1932), .IN3(n1955), .IN4(n973), .Q(g8774)
         );
  AO22X1 U2807 ( .IN1(g1633), .IN2(n1931), .IN3(n1955), .IN4(n970), .Q(g8777)
         );
  AO22X1 U2808 ( .IN1(g4), .IN2(n1975), .IN3(n1161), .IN4(n1162), .Q(g6656) );
  NOR2X0 U2809 ( .IN1(n1163), .IN2(n1164), .QN(n1162) );
  NOR4X0 U2810 ( .IN1(n1165), .IN2(n1707), .IN3(n1166), .IN4(n1628), .QN(n1161) );
  OR4X1 U2811 ( .IN1(g1466), .IN2(g1482), .IN3(g1486), .IN4(g1499), .Q(n1163)
         );
  AO22X1 U2812 ( .IN1(n650), .IN2(g682), .IN3(n1035), .IN4(g691), .Q(g8430) );
  AO22X1 U2813 ( .IN1(n624), .IN2(g1896), .IN3(n1039), .IN4(g1905), .Q(g8283)
         );
  AO22X1 U2814 ( .IN1(n650), .IN2(g691), .IN3(n1035), .IN4(g700), .Q(g8431) );
  AO22X1 U2815 ( .IN1(n624), .IN2(g1905), .IN3(n1039), .IN4(g1914), .Q(g8284)
         );
  AO22X1 U2816 ( .IN1(n650), .IN2(g664), .IN3(n1035), .IN4(g673), .Q(g8428) );
  AO22X1 U2817 ( .IN1(n624), .IN2(g1878), .IN3(n1039), .IN4(g1887), .Q(g8281)
         );
  AO22X1 U2818 ( .IN1(test_so7), .IN2(n1954), .IN3(g1027), .IN4(n1934), .Q(
        g6894) );
  AO22X1 U2819 ( .IN1(g1710), .IN2(n1954), .IN3(g1713), .IN4(n1933), .Q(g5396)
         );
  AO22X1 U2820 ( .IN1(g1080), .IN2(n1953), .IN3(g995), .IN4(n1936), .Q(g6895)
         );
  AO22X1 U2821 ( .IN1(g1083), .IN2(n1953), .IN3(g991), .IN4(n1934), .Q(g6898)
         );
  AO22X1 U2822 ( .IN1(g1089), .IN2(n1953), .IN3(test_so8), .IN4(n1935), .Q(
        g6908) );
  AO22X1 U2823 ( .IN1(g1086), .IN2(n1953), .IN3(g1003), .IN4(n1935), .Q(g6902)
         );
  AO22X1 U2824 ( .IN1(g1077), .IN2(n1953), .IN3(g1032), .IN4(n1938), .Q(g7257)
         );
  AO22X1 U2825 ( .IN1(g1071), .IN2(n1953), .IN3(g1023), .IN4(n1939), .Q(g7244)
         );
  AO22X1 U2826 ( .IN1(g1092), .IN2(n1953), .IN3(g1011), .IN4(n1938), .Q(g6912)
         );
  AO22X1 U2827 ( .IN1(g1074), .IN2(n1953), .IN3(g1015), .IN4(n1939), .Q(g6930)
         );
  AO22X1 U2828 ( .IN1(n1885), .IN2(n1953), .IN3(g1718), .IN4(n1937), .Q(g5404)
         );
  AO22X1 U2829 ( .IN1(g1095), .IN2(n1953), .IN3(test_so2), .IN4(n1936), .Q(
        g6918) );
  AO22X1 U2830 ( .IN1(g1098), .IN2(n1953), .IN3(g1019), .IN4(n1937), .Q(g6924)
         );
  AO22X1 U2831 ( .IN1(g1941), .IN2(n624), .IN3(n1039), .IN4(g1950), .Q(g8288)
         );
  AO22X1 U2832 ( .IN1(g727), .IN2(n650), .IN3(n1035), .IN4(g736), .Q(g8435) );
  AO21X1 U2833 ( .IN1(g1615), .IN2(n1958), .IN3(n565), .Q(n1067) );
  AO21X1 U2834 ( .IN1(g1621), .IN2(n1958), .IN3(n564), .Q(n1075) );
  AO21X1 U2835 ( .IN1(g1624), .IN2(n1959), .IN3(n563), .Q(n1080) );
  AO21X1 U2836 ( .IN1(g1639), .IN2(n1959), .IN3(n566), .Q(n1063) );
  AO21X1 U2837 ( .IN1(g1618), .IN2(n1958), .IN3(n567), .Q(n1084) );
  NAND3X0 U2838 ( .IN1(g611), .IN2(n1645), .IN3(g591), .QN(n805) );
  AO21X1 U2839 ( .IN1(g566), .IN2(n1958), .IN3(n568), .Q(g6035) );
  AO21X1 U2840 ( .IN1(g554), .IN2(n1958), .IN3(n566), .Q(g6000) );
  AO21X1 U2841 ( .IN1(g560), .IN2(n1958), .IN3(n564), .Q(g6015) );
  AO21X1 U2842 ( .IN1(g546), .IN2(n1958), .IN3(n567), .Q(g5996) );
  AO21X1 U2843 ( .IN1(g557), .IN2(n1958), .IN3(n565), .Q(g6002) );
  AO21X1 U2844 ( .IN1(g569), .IN2(n1958), .IN3(n569), .Q(g6038) );
  AO21X1 U2845 ( .IN1(g563), .IN2(n1958), .IN3(n563), .Q(g6026) );
  ISOLANDX1 U2846 ( .D(g4175), .ISO(n1214), .Q(n1193) );
  ISOLANDX1 U2847 ( .D(g4177), .ISO(n1153), .Q(n1125) );
  ISOLANDX1 U2848 ( .D(g4179), .ISO(n1099), .Q(n1093) );
  AO221X1 U2849 ( .IN1(g1878), .IN2(n1031), .IN3(g1950), .IN4(n624), .IN5(
        n1032), .Q(g8559) );
  AO221X1 U2850 ( .IN1(g664), .IN2(n1016), .IN3(g736), .IN4(n650), .IN5(n954), 
        .Q(g8649) );
  AO221X1 U2851 ( .IN1(n1104), .IN2(n959), .IN3(g639), .IN4(n649), .IN5(n954), 
        .Q(g7626) );
  NOR2X0 U2852 ( .IN1(g639), .IN2(n1105), .QN(n1104) );
  NOR4X0 U2853 ( .IN1(n719), .IN2(n720), .IN3(n834), .IN4(n717), .QN(n1105) );
  NAND2X0 U2854 ( .IN1(g682), .IN2(n899), .QN(n957) );
  NAND2X0 U2855 ( .IN1(g1896), .IN2(n853), .QN(n896) );
  NAND2X0 U2856 ( .IN1(g1905), .IN2(n853), .QN(n890) );
  NAND2X0 U2857 ( .IN1(g691), .IN2(n899), .QN(n948) );
  NAND3X0 U2858 ( .IN1(g374), .IN2(g369), .IN3(g378), .QN(n1385) );
  ISOLANDX1 U2859 ( .D(n1137), .ISO(g12), .Q(n1159) );
  ISOLANDX1 U2860 ( .D(g810), .ISO(n1151), .Q(n1123) );
  ISOLANDX1 U2861 ( .D(g818), .ISO(n1097), .Q(n1090) );
  XOR3X1 U2862 ( .IN1(n1869), .IN2(g1003), .IN3(n1870), .Q(n1398) );
  XNOR2X1 U2863 ( .IN1(g1015), .IN2(g1011), .Q(n1870) );
  NAND2X0 U2864 ( .IN1(g1700), .IN2(DFF_275_n1), .QN(g4089) );
  XOR3X1 U2865 ( .IN1(n1871), .IN2(g1019), .IN3(n1872), .Q(n1397) );
  XNOR2X1 U2866 ( .IN1(test_so8), .IN2(g995), .Q(n1872) );
  ISOLANDX1 U2867 ( .D(n817), .ISO(g1834), .Q(n1380) );
  NAND2X0 U2868 ( .IN1(n555), .IN2(g1766), .QN(n1175) );
  NAND2X0 U2869 ( .IN1(n1191), .IN2(g806), .QN(n1151) );
  NAND2X0 U2870 ( .IN1(n1123), .IN2(g814), .QN(n1097) );
  NOR2X0 U2871 ( .IN1(n1873), .IN2(n711), .QN(g4904) );
  NOR2X0 U2872 ( .IN1(n1874), .IN2(n667), .QN(g4892) );
  AND2X1 U2873 ( .IN1(g1703), .IN2(n560), .Q(n1875) );
  NAND3X0 U2874 ( .IN1(n906), .IN2(n908), .IN3(g722), .QN(n902) );
  NAND3X0 U2875 ( .IN1(n861), .IN2(n863), .IN3(g1936), .QN(n857) );
  NAND3X0 U2876 ( .IN1(n718), .IN2(n1693), .IN3(n907), .QN(n901) );
  NAND3X0 U2877 ( .IN1(n712), .IN2(n1694), .IN3(n862), .QN(n856) );
  AND4X1 U2878 ( .IN1(g658), .IN2(n934), .IN3(g668), .IN4(n967), .Q(n906) );
  ISOLANDX1 U2879 ( .D(g713), .ISO(n1656), .Q(n967) );
  AND4X1 U2880 ( .IN1(g1872), .IN2(n876), .IN3(g1882), .IN4(n921), .Q(n861) );
  ISOLANDX1 U2881 ( .D(g1927), .ISO(n1657), .Q(n921) );
  ISOLANDX1 U2882 ( .D(g1160), .ISO(n1967), .Q(g4334) );
  ISOLANDX1 U2883 ( .D(g1166), .ISO(n1967), .Q(g4325) );
  ISOLANDX1 U2884 ( .D(g148), .ISO(n1967), .Q(g6759) );
  ISOLANDX1 U2885 ( .D(g1157), .ISO(n1967), .Q(g4338) );
  ISOLANDX1 U2886 ( .D(g1163), .ISO(n1967), .Q(g4330) );
  ISOLANDX1 U2887 ( .D(g237), .ISO(n1967), .Q(g6821) );
  ISOLANDX1 U2888 ( .D(g1499), .ISO(n1967), .Q(g6198) );
  ISOLANDX1 U2889 ( .D(g1411), .ISO(n1967), .Q(g6244) );
  ISOLANDX1 U2890 ( .D(g225), .ISO(n1967), .Q(g6826) );
  ISOLANDX1 U2891 ( .D(g1407), .ISO(n1967), .Q(g6216) );
  ISOLANDX1 U2892 ( .D(g213), .ISO(n1966), .Q(g6829) );
  ISOLANDX1 U2893 ( .D(g186), .ISO(n1966), .Q(g6833) );
  ISOLANDX1 U2894 ( .D(g219), .ISO(n1966), .Q(g6827) );
  ISOLANDX1 U2895 ( .D(g143), .ISO(n1966), .Q(g6757) );
  ISOLANDX1 U2896 ( .D(g207), .ISO(n1966), .Q(g6831) );
  ISOLANDX1 U2897 ( .D(g231), .ISO(n1966), .Q(g6822) );
  ISOLANDX1 U2898 ( .D(g192), .ISO(n1966), .Q(g6838) );
  ISOLANDX1 U2899 ( .D(test_so3), .ISO(n1966), .Q(g6823) );
  ISOLANDX1 U2900 ( .D(g1371), .ISO(n1966), .Q(g6824) );
  ISOLANDX1 U2901 ( .D(g1383), .ISO(n1966), .Q(g6832) );
  ISOLANDX1 U2902 ( .D(g243), .ISO(n1966), .Q(g6819) );
  NOR2X0 U2903 ( .IN1(g1878), .IN2(n622), .QN(n922) );
  NOR2X0 U2904 ( .IN1(g664), .IN2(n648), .QN(n846) );
  AO21X1 U2905 ( .IN1(g119), .IN2(n1969), .IN3(n1195), .Q(g5918) );
  AO21X1 U2906 ( .IN1(g12), .IN2(n1969), .IN3(n1195), .Q(g5445) );
  AO21X1 U2907 ( .IN1(g9), .IN2(n1974), .IN3(n1195), .Q(g5421) );
  AO21X1 U2908 ( .IN1(n597), .IN2(n884), .IN3(n596), .Q(g8939) );
  XNOR2X1 U2909 ( .IN1(g1909), .IN2(n885), .Q(n884) );
  NAND2X0 U2910 ( .IN1(n855), .IN2(n886), .QN(n885) );
  AO222X1 U2911 ( .IN1(n875), .IN2(g1900), .IN3(n877), .IN4(n1675), .IN5(g1914), .IN6(n853), .Q(n886) );
  AO21X1 U2912 ( .IN1(n605), .IN2(n897), .IN3(n606), .Q(g8926) );
  XOR2X1 U2913 ( .IN1(g731), .IN2(n898), .Q(n897) );
  OA221X1 U2914 ( .IN1(g736), .IN2(n648), .IN3(n899), .IN4(n900), .IN5(n850), 
        .Q(n898) );
  NAND2X0 U2915 ( .IN1(n901), .IN2(n902), .QN(n900) );
  AO21X1 U2916 ( .IN1(n605), .IN2(n903), .IN3(n606), .Q(g8923) );
  XOR2X1 U2917 ( .IN1(g722), .IN2(n904), .Q(n903) );
  OA221X1 U2918 ( .IN1(g727), .IN2(n648), .IN3(n905), .IN4(n899), .IN5(n850), 
        .Q(n904) );
  OA22X1 U2919 ( .IN1(n718), .IN2(n906), .IN3(n907), .IN4(n908), .Q(n905) );
  AO21X1 U2920 ( .IN1(n597), .IN2(n851), .IN3(n596), .Q(g8945) );
  XOR2X1 U2921 ( .IN1(g1945), .IN2(n852), .Q(n851) );
  OA221X1 U2922 ( .IN1(g1950), .IN2(n622), .IN3(n853), .IN4(n854), .IN5(n855), 
        .Q(n852) );
  NAND2X0 U2923 ( .IN1(n856), .IN2(n857), .QN(n854) );
  AO21X1 U2924 ( .IN1(n597), .IN2(n858), .IN3(n596), .Q(g8944) );
  XOR2X1 U2925 ( .IN1(g1936), .IN2(n859), .Q(n858) );
  OA221X1 U2926 ( .IN1(g1941), .IN2(n622), .IN3(n860), .IN4(n853), .IN5(n855), 
        .Q(n859) );
  OA22X1 U2927 ( .IN1(n712), .IN2(n861), .IN3(n862), .IN4(n863), .Q(n860) );
  AO21X1 U2928 ( .IN1(n597), .IN2(n872), .IN3(n596), .Q(g8941) );
  XNOR2X1 U2929 ( .IN1(g1927), .IN2(n873), .Q(n872) );
  NAND2X0 U2930 ( .IN1(n855), .IN2(n874), .QN(n873) );
  AO222X1 U2931 ( .IN1(n875), .IN2(n876), .IN3(n877), .IN4(n878), .IN5(g1932), 
        .IN6(n853), .Q(n874) );
  AO21X1 U2932 ( .IN1(n1182), .IN2(n1029), .IN3(n1042), .Q(g6243) );
  OR2X1 U2933 ( .IN1(g798), .IN2(g794), .Q(n1182) );
  OA22X1 U2934 ( .IN1(g639), .IN2(n1024), .IN3(n1692), .IN4(n1025), .Q(n1023)
         );
  NOR3X0 U2935 ( .IN1(n1655), .IN2(g1840), .IN3(n1608), .QN(n809) );
  OR4X1 U2936 ( .IN1(g1240), .IN2(g1245), .IN3(g1235), .IN4(n1330), .Q(n1329)
         );
  OR3X1 U2937 ( .IN1(g1250), .IN2(g1260), .IN3(g1255), .Q(n1330) );
  OR4X1 U2938 ( .IN1(g391), .IN2(g396), .IN3(g386), .IN4(n1438), .Q(n1437) );
  OR3X1 U2939 ( .IN1(g401), .IN2(g411), .IN3(g406), .Q(n1438) );
  NAND2X0 U2940 ( .IN1(n1969), .IN2(n1058), .QN(n1040) );
  NAND3X0 U2941 ( .IN1(DFF_436_n1), .IN2(n594), .IN3(n1059), .QN(n1058) );
  NAND2X0 U2942 ( .IN1(n1969), .IN2(n1235), .QN(n1224) );
  NAND3X0 U2943 ( .IN1(n1236), .IN2(n1683), .IN3(g1212), .QN(n1235) );
  NAND2X0 U2944 ( .IN1(n1090), .IN2(g822), .QN(n1043) );
  NBUFFX2 U2945 ( .IN(g1713), .Q(n1885) );
  NAND2X0 U2946 ( .IN1(n520), .IN2(g794), .QN(g5849) );
  NAND3X0 U2947 ( .IN1(n804), .IN2(g605), .IN3(n721), .QN(n837) );
  AOI22X1 U2948 ( .IN1(n1876), .IN2(n1877), .IN3(n1878), .IN4(g431), .QN(n1434) );
  OAI21X1 U2949 ( .IN1(n1436), .IN2(n1437), .IN3(n1878), .QN(n1877) );
  OA21X1 U2950 ( .IN1(n1052), .IN2(n1053), .IN3(n1610), .Q(g8173) );
  OA21X1 U2951 ( .IN1(n1054), .IN2(n1055), .IN3(g1806), .Q(n1053) );
  AND3X1 U2952 ( .IN1(n1056), .IN2(n1055), .IN3(g1801), .Q(n1052) );
  NAND3X0 U2953 ( .IN1(g1801), .IN2(n1057), .IN3(g1806), .QN(n1055) );
  OR4X1 U2954 ( .IN1(test_so6), .IN2(g1275), .IN3(g1265), .IN4(n1331), .Q(
        n1328) );
  OR4X1 U2955 ( .IN1(g1304), .IN2(g1300), .IN3(g1296), .IN4(g1292), .Q(n1331)
         );
  OR4X1 U2956 ( .IN1(g421), .IN2(g426), .IN3(g416), .IN4(n1439), .Q(n1436) );
  OR4X1 U2957 ( .IN1(g452), .IN2(g448), .IN3(g444), .IN4(g440), .Q(n1439) );
  NOR2X0 U2958 ( .IN1(n1041), .IN2(n1042), .QN(g8245) );
  XOR2X1 U2959 ( .IN1(n1043), .IN2(g826), .Q(n1041) );
  OAI22X1 U2960 ( .IN1(g525), .IN2(n1698), .IN3(g521), .IN4(n1354), .QN(n1241)
         );
  OA21X1 U2961 ( .IN1(n1355), .IN2(n1356), .IN3(n1695), .Q(n1354) );
  NOR2X0 U2962 ( .IN1(n954), .IN2(n961), .QN(g8820) );
  XOR2X1 U2963 ( .IN1(n603), .IN2(g622), .Q(n961) );
  NAND3X0 U2964 ( .IN1(g4892), .IN2(n1020), .IN3(n1021), .QN(n1019) );
  NAND4X0 U2965 ( .IN1(n1024), .IN2(n1026), .IN3(n953), .IN4(n1025), .QN(n1020) );
  XOR2X1 U2966 ( .IN1(n1022), .IN2(n1023), .Q(n1021) );
  NAND2X0 U2967 ( .IN1(g255), .IN2(g622), .QN(n1022) );
  NAND3X0 U2968 ( .IN1(n1118), .IN2(n1119), .IN3(n643), .QN(g7441) );
  NAND2X0 U2969 ( .IN1(g643), .IN2(n1701), .QN(n1118) );
  INVX0 U2970 ( .IN(n1101), .QN(n643) );
  NOR2X0 U2971 ( .IN1(n1964), .IN2(n1062), .QN(g8055) );
  XNOR2X1 U2972 ( .IN1(g1490), .IN2(n1063), .Q(n1062) );
  NOR2X0 U2973 ( .IN1(n1963), .IN2(n1078), .QN(g8044) );
  XNOR2X1 U2974 ( .IN1(g131), .IN2(g6038), .Q(n1078) );
  NOR2X0 U2975 ( .IN1(n1964), .IN2(n1064), .QN(g8054) );
  XNOR2X1 U2976 ( .IN1(g174), .IN2(g6015), .Q(n1064) );
  NOR2X0 U2977 ( .IN1(n1983), .IN2(n1065), .QN(g8053) );
  XNOR2X1 U2978 ( .IN1(g139), .IN2(g6045), .Q(n1065) );
  NOR2X0 U2979 ( .IN1(n1964), .IN2(n1061), .QN(g8059) );
  XNOR2X1 U2980 ( .IN1(g135), .IN2(g6042), .Q(n1061) );
  NOR2X0 U2981 ( .IN1(n1983), .IN2(n1066), .QN(g8052) );
  XNOR2X1 U2982 ( .IN1(g1486), .IN2(n1067), .Q(n1066) );
  NOR2X0 U2983 ( .IN1(n1966), .IN2(n1071), .QN(g8049) );
  XNOR2X1 U2984 ( .IN1(g166), .IN2(g6049), .Q(n1071) );
  NOR2X0 U2985 ( .IN1(n1983), .IN2(n1072), .QN(g8048) );
  XNOR2X1 U2986 ( .IN1(g153), .IN2(g5996), .Q(n1072) );
  NOR2X0 U2987 ( .IN1(n1962), .IN2(n1079), .QN(g8043) );
  XNOR2X1 U2988 ( .IN1(g1478), .IN2(n1080), .Q(n1079) );
  NOR2X0 U2989 ( .IN1(n1962), .IN2(n1085), .QN(g8040) );
  XNOR2X1 U2990 ( .IN1(g1474), .IN2(n1086), .Q(n1085) );
  NOR2X0 U2991 ( .IN1(n1963), .IN2(n972), .QN(g8775) );
  XNOR2X1 U2992 ( .IN1(g1436), .IN2(n973), .Q(n972) );
  NOR2X0 U2993 ( .IN1(n1964), .IN2(n1060), .QN(g8060) );
  XNOR2X1 U2994 ( .IN1(g162), .IN2(g6002), .Q(n1060) );
  NOR2X0 U2995 ( .IN1(n1962), .IN2(n1087), .QN(g8039) );
  XNOR2X1 U2996 ( .IN1(g1470), .IN2(n1088), .Q(n1087) );
  NOR2X0 U2997 ( .IN1(n1962), .IN2(n1095), .QN(g7843) );
  XNOR2X1 U2998 ( .IN1(g158), .IN2(g6000), .Q(n1095) );
  NOR2X0 U2999 ( .IN1(n1962), .IN2(n1076), .QN(g8045) );
  XNOR2X1 U3000 ( .IN1(g1462), .IN2(n1077), .Q(n1076) );
  NOR2X0 U3001 ( .IN1(n1962), .IN2(n988), .QN(g8769) );
  XNOR2X1 U3002 ( .IN1(g1428), .IN2(n987), .Q(n988) );
  NOR2X0 U3003 ( .IN1(n1983), .IN2(n1070), .QN(g8050) );
  XNOR2X1 U3004 ( .IN1(g170), .IN2(g6026), .Q(n1070) );
  NOR2X0 U3005 ( .IN1(n1983), .IN2(n1068), .QN(g8051) );
  XNOR2X1 U3006 ( .IN1(g1466), .IN2(n1069), .Q(n1068) );
  NOR2X0 U3007 ( .IN1(n1962), .IN2(n1074), .QN(g8046) );
  XNOR2X1 U3008 ( .IN1(g1482), .IN2(n1075), .Q(n1074) );
  NOR2X0 U3009 ( .IN1(n1966), .IN2(n1006), .QN(g8766) );
  XNOR2X1 U3010 ( .IN1(g1448), .IN2(n969), .Q(n1006) );
  NOR2X0 U3011 ( .IN1(n1962), .IN2(n1083), .QN(g8041) );
  XNOR2X1 U3012 ( .IN1(g1494), .IN2(n1084), .Q(n1083) );
  NBUFFX2 U3013 ( .IN(g1690), .Q(n1882) );
  NOR2X0 U3014 ( .IN1(n1961), .IN2(n994), .QN(g8768) );
  XNOR2X1 U3015 ( .IN1(g1444), .IN2(n970), .Q(n994) );
  NOR2X0 U3016 ( .IN1(n1961), .IN2(n1011), .QN(g8765) );
  XNOR2X1 U3017 ( .IN1(g1432), .IN2(n979), .Q(n1011) );
  NOR2X0 U3018 ( .IN1(n1961), .IN2(n1000), .QN(g8767) );
  XNOR2X1 U3019 ( .IN1(g1403), .IN2(n986), .Q(n1000) );
  NOR2X0 U3020 ( .IN1(n1961), .IN2(n980), .QN(g8772) );
  XNOR2X1 U3021 ( .IN1(g1440), .IN2(n971), .Q(n980) );
  NOR4X0 U3022 ( .IN1(n1275), .IN2(n1276), .IN3(n1277), .IN4(n1278), .QN(n1274) );
  XOR2X1 U3023 ( .IN1(test_so8), .IN2(g1245), .Q(n1276) );
  XOR2X1 U3024 ( .IN1(g991), .IN2(g1235), .Q(n1278) );
  XOR2X1 U3025 ( .IN1(g1250), .IN2(g1011), .Q(n1277) );
  NOR4X0 U3026 ( .IN1(n1425), .IN2(n1426), .IN3(n1427), .IN4(n1428), .QN(n1424) );
  XOR2X1 U3027 ( .IN1(g396), .IN2(g324), .Q(n1426) );
  XOR2X1 U3028 ( .IN1(g386), .IN2(g318), .Q(n1428) );
  XOR2X1 U3029 ( .IN1(g401), .IN2(g327), .Q(n1427) );
  NOR4X0 U3030 ( .IN1(g1166), .IN2(g1163), .IN3(g1160), .IN4(g1157), .QN(n1269) );
  NBUFFX2 U3031 ( .IN(g456), .Q(n1884) );
  NOR3X0 U3032 ( .IN1(g1909), .IN2(g1918), .IN3(g1900), .QN(n878) );
  NOR3X0 U3033 ( .IN1(g695), .IN2(g704), .IN3(g686), .QN(n936) );
  NOR3X0 U3034 ( .IN1(g1861), .IN2(g1864), .IN3(n1642), .QN(n1147) );
  NOR2X0 U3035 ( .IN1(n711), .IN2(DFF_489_n1), .QN(g4905) );
  NOR2X0 U3036 ( .IN1(n711), .IN2(DFF_385_n1), .QN(g4902) );
  NOR2X0 U3037 ( .IN1(n711), .IN2(DFF_330_n1), .QN(g4903) );
  NOR2X0 U3038 ( .IN1(n667), .IN2(DFF_157_n1), .QN(g4893) );
  NOR2X0 U3039 ( .IN1(n667), .IN2(DFF_336_n1), .QN(g4890) );
  NOR2X0 U3040 ( .IN1(n667), .IN2(DFF_136_n1), .QN(g4891) );
  NOR2X0 U3041 ( .IN1(n1199), .IN2(n1961), .QN(g5755) );
  XOR3X1 U3042 ( .IN1(g1389), .IN2(n1200), .IN3(n1201), .Q(n1199) );
  XOR2X1 U3043 ( .IN1(g201), .IN2(g197), .Q(n1201) );
  NOR2X0 U3044 ( .IN1(g1386), .IN2(n1202), .QN(n1200) );
  NOR2X0 U3045 ( .IN1(n1179), .IN2(n1961), .QN(g6439) );
  XNOR3X1 U3046 ( .IN1(n1180), .IN2(g153), .IN3(g182), .Q(n1179) );
  XOR2X1 U3047 ( .IN1(g148), .IN2(g143), .Q(n1180) );
  NOR2X0 U3048 ( .IN1(n1196), .IN2(n1961), .QN(g5770) );
  XOR3X1 U3049 ( .IN1(n1197), .IN2(g1499), .IN3(n1707), .Q(n1196) );
  XOR2X1 U3050 ( .IN1(g1494), .IN2(g1453), .Q(n1197) );
  OR2X1 U3051 ( .IN1(g1900), .IN2(g1909), .Q(n882) );
  OR2X1 U3052 ( .IN1(g686), .IN2(g695), .Q(n940) );
  NAND2X0 U3053 ( .IN1(n995), .IN2(n996), .QN(n970) );
  AO221X1 U3054 ( .IN1(n997), .IN2(g1141), .IN3(n1660), .IN4(n998), .IN5(g2355), .Q(n996) );
  NOR2X0 U3055 ( .IN1(g1101), .IN2(n999), .QN(n997) );
  NAND2X0 U3056 ( .IN1(n634), .IN2(n1654), .QN(n998) );
  NAND2X0 U3057 ( .IN1(n981), .IN2(n982), .QN(n971) );
  AO221X1 U3058 ( .IN1(n983), .IN2(g1137), .IN3(n1597), .IN4(n984), .IN5(g2355), .Q(n982) );
  NAND2X0 U3059 ( .IN1(n631), .IN2(g1101), .QN(n984) );
  NOR2X0 U3060 ( .IN1(n1654), .IN2(n978), .QN(n983) );
  NAND2X0 U3061 ( .IN1(n989), .IN2(n990), .QN(n987) );
  AO221X1 U3062 ( .IN1(n991), .IN2(g1121), .IN3(n1618), .IN4(n992), .IN5(g2355), .Q(n990) );
  NOR2X0 U3063 ( .IN1(n1654), .IN2(n993), .QN(n991) );
  NAND2X0 U3064 ( .IN1(n632), .IN2(g1101), .QN(n992) );
  AND4X1 U3065 ( .IN1(n1625), .IN2(n1688), .IN3(n1208), .IN4(n1209), .Q(n1184)
         );
  NOR2X0 U3066 ( .IN1(g1371), .IN2(test_so3), .QN(n1208) );
  NOR4X0 U3067 ( .IN1(g243), .IN2(g237), .IN3(g231), .IN4(g225), .QN(n1209) );
  AO21X1 U3068 ( .IN1(n605), .IN2(n942), .IN3(n606), .Q(g8887) );
  XNOR2X1 U3069 ( .IN1(g695), .IN2(n943), .Q(n942) );
  NAND2X0 U3070 ( .IN1(n850), .IN2(n944), .QN(n943) );
  AO222X1 U3071 ( .IN1(n933), .IN2(g686), .IN3(n935), .IN4(n1676), .IN5(g700), 
        .IN6(n899), .Q(n944) );
  NOR2X0 U3072 ( .IN1(n1191), .IN2(n1212), .QN(g5543) );
  OA22X1 U3073 ( .IN1(n1622), .IN2(n1042), .IN3(g5849), .IN4(n1717), .Q(n1212)
         );
  XNOR2X1 U3074 ( .IN1(test_so1), .IN2(n1045), .Q(N599) );
  NOR3X0 U3075 ( .IN1(g1125), .IN2(g1133), .IN3(g1129), .QN(n1268) );
  AO21X1 U3076 ( .IN1(n597), .IN2(n879), .IN3(n596), .Q(g8940) );
  XOR2X1 U3077 ( .IN1(g1918), .IN2(n880), .Q(n879) );
  NOR2X0 U3078 ( .IN1(n881), .IN2(n620), .QN(n880) );
  OA222X1 U3079 ( .IN1(n622), .IN2(n1718), .IN3(n600), .IN4(n882), .IN5(n595), 
        .IN6(n883), .Q(n881) );
  AO21X1 U3080 ( .IN1(n605), .IN2(n937), .IN3(n606), .Q(g8889) );
  XOR2X1 U3081 ( .IN1(g704), .IN2(n938), .Q(n937) );
  NOR2X0 U3082 ( .IN1(n939), .IN2(n644), .QN(n938) );
  OA222X1 U3083 ( .IN1(n648), .IN2(n1719), .IN3(n645), .IN4(n940), .IN5(n646), 
        .IN6(n941), .Q(n939) );
  NOR3X0 U3084 ( .IN1(n1431), .IN2(n1432), .IN3(n1433), .QN(n1423) );
  XOR2X1 U3085 ( .IN1(g421), .IN2(g312), .Q(n1431) );
  XOR2X1 U3086 ( .IN1(g411), .IN2(g333), .Q(n1433) );
  XOR2X1 U3087 ( .IN1(n1681), .IN2(n1390), .Q(n1432) );
  NBUFFX2 U3088 ( .IN(g456), .Q(n1883) );
  NOR3X0 U3089 ( .IN1(n1150), .IN2(n1123), .IN3(n1042), .QN(g6733) );
  ISOLANDX1 U3090 ( .D(n1151), .ISO(g810), .Q(n1150) );
  NOR3X0 U3091 ( .IN1(n1096), .IN2(n1090), .IN3(n1042), .QN(g7709) );
  ISOLANDX1 U3092 ( .D(n1097), .ISO(g818), .Q(n1096) );
  NOR3X0 U3093 ( .IN1(n1098), .IN2(n1093), .IN3(n537), .QN(g7705) );
  ISOLANDX1 U3094 ( .D(n1099), .ISO(g4179), .Q(n1098) );
  NOR3X0 U3095 ( .IN1(n1213), .IN2(n1193), .IN3(n537), .QN(g5536) );
  ISOLANDX1 U3096 ( .D(n1214), .ISO(g4175), .Q(n1213) );
  NOR3X0 U3097 ( .IN1(n1152), .IN2(n1125), .IN3(n537), .QN(g6728) );
  ISOLANDX1 U3098 ( .D(n1153), .ISO(g4177), .Q(n1152) );
  NAND4X0 U3099 ( .IN1(n1159), .IN2(g1470), .IN3(g1474), .IN4(g1494), .QN(
        n1165) );
  NBUFFX2 U3100 ( .IN(g1690), .Q(n1881) );
  NOR2X0 U3101 ( .IN1(n1885), .IN2(n1174), .QN(g6508) );
  OA22X1 U3102 ( .IN1(n1175), .IN2(n1176), .IN3(n553), .IN4(n1715), .Q(n1174)
         );
  NAND2X0 U3103 ( .IN1(test_so5), .IN2(n1172), .QN(n1176) );
  NOR2X0 U3104 ( .IN1(n1885), .IN2(n1138), .QN(g6983) );
  OA22X1 U3105 ( .IN1(n1139), .IN2(n1140), .IN3(n1116), .IN4(n1702), .Q(n1138)
         );
  NAND2X0 U3106 ( .IN1(g1786), .IN2(n1117), .QN(n1140) );
  NAND4X0 U3107 ( .IN1(n1679), .IN2(n1620), .IN3(n1600), .IN4(n1358), .QN(
        n1355) );
  NOR4X0 U3108 ( .IN1(g542), .IN2(g538), .IN3(g534), .IN4(g530), .QN(n1358) );
  NOR2X0 U3109 ( .IN1(n1885), .IN2(n1094), .QN(g7930) );
  XNOR2X1 U3110 ( .IN1(n1056), .IN2(g1801), .Q(n1094) );
  NOR2X0 U3111 ( .IN1(n1957), .IN2(n818), .QN(g9269) );
  XOR2X1 U3112 ( .IN1(g1822), .IN2(n819), .Q(n818) );
  NOR2X0 U3113 ( .IN1(n820), .IN2(n821), .QN(n819) );
  AOI21X1 U3114 ( .IN1(n822), .IN2(n815), .IN3(n598), .QN(n821) );
  NOR2X0 U3115 ( .IN1(n1958), .IN2(n1033), .QN(g8505) );
  XOR2X1 U3116 ( .IN1(g617), .IN2(n1034), .Q(n1033) );
  AOI21X1 U3117 ( .IN1(n650), .IN2(g736), .IN3(n960), .QN(n1034) );
  NOR2X0 U3118 ( .IN1(n1958), .IN2(n800), .QN(g9721) );
  XOR2X1 U3119 ( .IN1(g611), .IN2(n801), .Q(n800) );
  OA21X1 U3120 ( .IN1(n802), .IN2(n649), .IN3(n803), .Q(n801) );
  OA21X1 U3121 ( .IN1(n804), .IN2(n805), .IN3(n1645), .Q(n802) );
  NOR2X0 U3122 ( .IN1(n1957), .IN2(n835), .QN(g9124) );
  XOR2X1 U3123 ( .IN1(g599), .IN2(n836), .Q(n835) );
  ISOLANDX1 U3124 ( .D(n837), .ISO(n838), .Q(n836) );
  OA21X1 U3125 ( .IN1(n720), .IN2(n717), .IN3(n804), .Q(n838) );
  NOR2X0 U3126 ( .IN1(n1957), .IN2(n823), .QN(g9266) );
  XOR2X1 U3127 ( .IN1(g1814), .IN2(n824), .Q(n823) );
  NOR2X0 U3128 ( .IN1(n825), .IN2(n820), .QN(n824) );
  OA21X1 U3129 ( .IN1(n809), .IN2(n713), .IN3(n812), .Q(n825) );
  NOR2X0 U3130 ( .IN1(n1885), .IN2(n1177), .QN(g6502) );
  XOR2X1 U3131 ( .IN1(n1175), .IN2(test_so5), .Q(n1177) );
  NOR2X0 U3132 ( .IN1(n1885), .IN2(n1168), .QN(g6525) );
  XOR2X1 U3133 ( .IN1(n1139), .IN2(g1786), .Q(n1168) );
  NOR2X0 U3134 ( .IN1(n1958), .IN2(n1036), .QN(g8384) );
  XOR2X1 U3135 ( .IN1(g1840), .IN2(n1037), .Q(n1036) );
  AOI21X1 U3136 ( .IN1(n624), .IN2(g1950), .IN3(n929), .QN(n1037) );
  NAND4X0 U3137 ( .IN1(n1680), .IN2(n1621), .IN3(n1599), .IN4(n1357), .QN(
        n1356) );
  NOR3X0 U3138 ( .IN1(g491), .IN2(g501), .IN3(g496), .QN(n1357) );
  INVX0 U3139 ( .IN(g23), .QN(g3327) );
  INVX0 U3140 ( .IN(g18), .QN(n1960) );
  NAND2X0 U3141 ( .IN1(n1279), .IN2(n1280), .QN(n1275) );
  XNOR2X1 U3142 ( .IN1(g995), .IN2(g1275), .Q(n1279) );
  XNOR2X1 U3143 ( .IN1(g1003), .IN2(g1240), .Q(n1280) );
  NAND2X0 U3144 ( .IN1(n1429), .IN2(n1430), .QN(n1425) );
  XNOR2X1 U3145 ( .IN1(g315), .IN2(g426), .Q(n1429) );
  XNOR2X1 U3146 ( .IN1(g321), .IN2(g391), .Q(n1430) );
  INVX0 U3147 ( .IN(g881), .QN(n594) );
  NAND2X0 U3148 ( .IN1(g1703), .IN2(n1724), .QN(n1451) );
  NAND2X0 U3149 ( .IN1(n1229), .IN2(g1351), .QN(n1228) );
  NAND2X0 U3150 ( .IN1(n617), .IN2(g986), .QN(n1338) );
  AND3X1 U3151 ( .IN1(g1336), .IN2(g1346), .IN3(g1341), .Q(n1229) );
  NAND3X0 U3152 ( .IN1(n1612), .IN2(n1595), .IN3(g650), .QN(n1129) );
  NAND3X0 U3153 ( .IN1(g971), .IN2(g981), .IN3(g976), .QN(n1342) );
  NAND2X0 U3154 ( .IN1(g1909), .IN2(g1900), .QN(n883) );
  NAND2X0 U3155 ( .IN1(g695), .IN2(g686), .QN(n941) );
  AO22X1 U3156 ( .IN1(g1786), .IN2(n725), .IN3(g1750), .IN4(n1217), .Q(g4264)
         );
  AO22X1 U3157 ( .IN1(g1796), .IN2(n725), .IN3(g1756), .IN4(n1217), .Q(g4283)
         );
  AO22X1 U3158 ( .IN1(g1781), .IN2(n725), .IN3(g1747), .IN4(n1217), .Q(g4255)
         );
  AO22X1 U3159 ( .IN1(g1806), .IN2(n725), .IN3(g1762), .IN4(n1217), .Q(g4309)
         );
  AO22X1 U3160 ( .IN1(g1766), .IN2(n725), .IN3(g1738), .IN4(n1217), .Q(g4231)
         );
  AO22X1 U3161 ( .IN1(g1791), .IN2(n725), .IN3(g1753), .IN4(n1217), .Q(g4274)
         );
  AO22X1 U3162 ( .IN1(test_so5), .IN2(n725), .IN3(g1741), .IN4(n1217), .Q(
        g4238) );
  AO22X1 U3163 ( .IN1(g1801), .IN2(n725), .IN3(g1759), .IN4(n1217), .Q(g4293)
         );
  AO22X1 U3164 ( .IN1(g1776), .IN2(n725), .IN3(g1744), .IN4(n1217), .Q(g4239)
         );
  NAND4X0 U3165 ( .IN1(g1444), .IN2(g1428), .IN3(g1440), .IN4(g1436), .QN(
        n1157) );
  NAND4X0 U3166 ( .IN1(g1478), .IN2(g1462), .IN3(g1490), .IN4(n1703), .QN(
        n1164) );
  NAND2X0 U3167 ( .IN1(g806), .IN2(g802), .QN(n1030) );
  NOR2X0 U3168 ( .IN1(g1737), .IN2(g1610), .QN(g2478) );
  NOR2X0 U3169 ( .IN1(n562), .IN2(n1189), .QN(g6155) );
  XOR2X1 U3170 ( .IN1(g1707), .IN2(n1653), .Q(n1189) );
  ISOLANDX1 U3171 ( .D(g1610), .ISO(n555), .Q(g5194) );
  NAND2X0 U3172 ( .IN1(n1131), .IN2(n1610), .QN(g7133) );
  XOR2X1 U3173 ( .IN1(g1766), .IN2(n1054), .Q(n1131) );
  AO21X1 U3174 ( .IN1(g654), .IN2(n1100), .IN3(n1101), .Q(g7660) );
  NAND4X0 U3175 ( .IN1(g627), .IN2(n1612), .IN3(n1595), .IN4(n1709), .QN(n1100) );
  AO21X1 U3176 ( .IN1(g1868), .IN2(n1143), .IN3(n1144), .Q(g6909) );
  OR3X1 U3177 ( .IN1(g1861), .IN2(g1864), .IN3(n1642), .Q(n1143) );
  OA21X1 U3178 ( .IN1(n1146), .IN2(n1147), .IN3(n619), .Q(g6795) );
  OA21X1 U3179 ( .IN1(g1861), .IN2(n1642), .IN3(g1864), .Q(n1146) );
  OA21X1 U3180 ( .IN1(n1218), .IN2(n592), .IN3(g746), .Q(g3462) );
  NOR2X0 U3181 ( .IN1(g750), .IN2(n1647), .QN(n1218) );
  NOR2X0 U3182 ( .IN1(n1178), .IN2(n1144), .QN(g6471) );
  XOR2X1 U3183 ( .IN1(n1642), .IN2(g1861), .Q(n1178) );
  NOR4X0 U3184 ( .IN1(n1210), .IN2(n1211), .IN3(n1702), .IN4(n1626), .QN(g5556) );
  NAND4X0 U3185 ( .IN1(n1882), .IN2(g1707), .IN3(g1806), .IN4(g1801), .QN(
        n1210) );
  NAND3X0 U3186 ( .IN1(n661), .IN2(n1659), .IN3(g1786), .QN(n1211) );
  NOR2X0 U3187 ( .IN1(g1707), .IN2(n562), .QN(g4076) );
  NAND2X0 U3188 ( .IN1(g814), .IN2(g810), .QN(n1028) );
  NAND2X0 U3189 ( .IN1(g822), .IN2(g818), .QN(n1027) );
  NAND4X0 U3190 ( .IN1(g170), .IN2(g174), .IN3(n1613), .IN4(n1704), .QN(n1135)
         );
  OR2X1 U3191 ( .IN1(g1289), .IN2(g1212), .Q(g4556) );
  INVX0 U3192 ( .IN(g1700), .QN(n562) );

  // Trojan trigger ----------------
  AND2X2 Tg1_Trojan1 (.IN1(g6179), .IN2(n519), .Q(Tg1_OUT1));
  AND2X2 Tg1_Trojan2 (.IN1(n1202), .IN2(n1132), .Q(Tg1_OUT2));
  AND2X2 Tg1_Trojan3 (.IN1(n1226), .IN2(n1858), .Q(Tg1_OUT3));
  AND2X2 Tg1_Trojan4 (.IN1(g5556), .IN2(n898), .Q(Tg1_OUT4));
  AND4X1 Tg1_Trojan1234 (.IN1(Tg1_OUT1), .IN2(Tg1_OUT2), .IN3(Tg1_OUT3), .IN4(Tg1_OUT4), .Q(Tg1_OUT1234));
  NOR2X0 Tg1_Trojan5 (.IN1(n1391), .IN2(n931), .QN(Tg1_OUT5));
  NOR2X0 Tg1_Trojan6 (.IN1(n857), .IN2(n902), .QN(Tg1_OUT6));
  NOR2X0 Tg1_Trojan7 (.IN1(n1889), .IN2(n1890), .QN(Tg1_OUT7));
  NOR2X0 Tg1_Trojan8 (.IN1(n1055), .IN2(n1016), .QN(Tg1_OUT8));
  AND4X1 Tg1_Trojan5678 (.IN1(Tg1_OUT5), .IN2(Tg1_OUT6), .IN3(Tg1_OUT7), .IN4(Tg1_OUT8), .Q(Tg1_OUT5678));
  AND2X2 Tg1_Tj_Trigger ( .IN1(Tg1_OUT1234), .IN2(Tg1_OUT5678), .Q(Tg1_Trigger1) );
  DFFNX2 Tg1_Trigger ( .CLK(Tg1_Trigger1), .D(1'b1), .Q(Tg1) ); 

  AND2X2 Tg2_Trojan1 (.IN1(n938), .IN2(n1917), .Q(Tg2_OUT1));
  AND2X2 Tg2_Trojan2 (.IN1(n1921), .IN2(n1911), .Q(Tg2_OUT2));
  AND2X2 Tg2_Trojan3 (.IN1(n1918), .IN2(n1913), .Q(Tg2_OUT3));
  AND2X2 Tg2_Trojan4 (.IN1(n1916), .IN2(n1910), .Q(Tg2_OUT4));
  AND4X1 Tg2_Trojan1234 (.IN1(Tg2_OUT1), .IN2(Tg2_OUT2), .IN3(Tg2_OUT3), .IN4(Tg2_OUT4), .Q(Tg2_OUT1234));
  AND2X2 Tg2_Trojan5 (.IN1(n1161), .IN2(n1154), .Q(Tg2_OUT5));
  AND2X2 Tg2_Trojan6 (.IN1(n1116), .IN2(n1162), .Q(Tg2_OUT6));
  AND2X2 Tg2_Trojan7 (.IN1(n1155), .IN2(n1107), .Q(Tg2_OUT7));
  AND2X2 Tg2_Trojan8 (.IN1(n929), .IN2(n554), .Q(Tg2_OUT8));
  AND4X1 Tg2_Trojan5678 (.IN1(Tg2_OUT5), .IN2(Tg2_OUT6), .IN3(Tg2_OUT7), .IN4(Tg2_OUT8), .Q(Tg2_OUT5678));
  AND2X2 Tg2_Tj_Trigger ( .IN1(Tg2_OUT1234), .IN2(Tg2_OUT5678), .Q(Tg2_Trigger2) );
  DFFNX2 Tg2_Trigger ( .CLK(Tg2_Trigger2), .D(Tg1), .Q(Tg2) ); 

  INVX0 INVtest_se ( .IN(test_se), .QN(test_se_NOT) );
  AND2X2 Trojan_Trigger (.IN1(Tg2), .IN2(test_se_NOT), .Q(Trigger_select) );

  // Trojan payload ----------------
  MUX21X2 Trojan_Paylaod ( .IN1(g4207_Payload), .IN2(n1936), .S(Trigger_select), .Q(g4207) );

endmodule

